----------------------------------------------------------
--
-- 32 bits pipelined RISC processor
-- Copyright (c) 2010 Victor Munoz. All rights reserved.
-- derechos reservados, prohibida su reproduccion
--
-- Author: Victor Munoz
-- Contact: vmunoz@ingenieria-inversa.cl
--
----------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

----------------------------------------------------------

ENTITY SRAM IS
    GENERIC(
        ADDR:     INTEGER:= (9+2);
        DEPTH:    INTEGER:= 512
    );
    PORT(
        CLK:      IN  STD_LOGIC;
        ENABLE:   IN  STD_LOGIC;
        R:        IN  STD_LOGIC;
        W:        IN  STD_LOGIC;
        RADDR:    IN  STD_LOGIC_VECTOR(ADDR-1 DOWNTO 0);
        WADDR:    IN  STD_LOGIC_VECTOR(ADDR-1 DOWNTO 0);
        DATA_IN:  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
        MODE:     IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
        ISSIGNED: IN  STD_LOGIC;
        DATA_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0):= "00000000000000000000000000000000"
    );
END SRAM;

--------------------------------------------------------------

ARCHITECTURE BEHAV_CODE OF SRAM IS

    TYPE RAM_TYPE IS ARRAY (0 TO DEPTH-1) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL TMP_RAM: RAM_TYPE := (

         0 => x"3C080000", -- lui $t0, 0000
         1 => x"2508084C", -- addiu $t0, $t0, 2124
         2 => x"3C090000", -- lui $t1, 0000
         3 => x"25290854", -- addiu $t1, $t1, 2132
         4 => x"11090003", -- beq $t0, $t1, 3
         5 => x"25080004", -- addiu $t0, $t0, 4
         6 => x"08000004", -- j 4
         7 => x"AD00FFFC", -- sw $zero, -4(t0)
         8 => x"00000821", -- addu $at, $zero, $zero
         9 => x"00001021", -- addu $v0, $zero, $zero
        10 => x"00001821", -- addu $v1, $zero, $zero
        11 => x"00002021", -- addu $a0, $zero, $zero
        12 => x"00002821", -- addu $a1, $zero, $zero
        13 => x"00003021", -- addu $a2, $zero, $zero
        14 => x"00003821", -- addu $a3, $zero, $zero
        15 => x"00004021", -- addu $t0, $zero, $zero
        16 => x"00004821", -- addu $t1, $zero, $zero
        17 => x"00005021", -- addu $t2, $zero, $zero
        18 => x"00005821", -- addu $t3, $zero, $zero
        19 => x"00006021", -- addu $t4, $zero, $zero
        20 => x"00006821", -- addu $t5, $zero, $zero
        21 => x"00007021", -- addu $t6, $zero, $zero
        22 => x"00007821", -- addu $t7, $zero, $zero
        23 => x"00008021", -- addu $s0, $zero, $zero
        24 => x"00008821", -- addu $s1, $zero, $zero
        25 => x"00009021", -- addu $s2, $zero, $zero
        26 => x"00009821", -- addu $s3, $zero, $zero
        27 => x"0000A021", -- addu $s4, $zero, $zero
        28 => x"0000A821", -- addu $s5, $zero, $zero
        29 => x"0000B021", -- addu $s6, $zero, $zero
        30 => x"0000B821", -- addu $s7, $zero, $zero
        31 => x"0000C021", -- addu $t8, $zero, $zero
        32 => x"0000C821", -- addu $t9, $zero, $zero
        33 => x"0000D021", -- addu $k0, $zero, $zero
        34 => x"0000D821", -- addu $k1, $zero, $zero
        35 => x"0000E021", -- addu $gp, $zero, $zero
        36 => x"0000F821", -- addu $ra, $zero, $zero
        37 => x"3C1D0000", -- lui $sp, 0000
        38 => x"27BD0FF8", -- addiu $sp, $sp, 4088
        39 => x"0C0001CD", -- jal 461
        40 => x"03A0F021", -- addu $fp, $sp, $zero
        41 => x"08000029", -- j 41
        42 => x"00000000", -- nop
        43 => x"27BDFFF8", -- addiu $sp, $sp, -8
        44 => x"AFBE0004", -- sw $fp, 4(sp)
        45 => x"03A0F021", -- addu $fp, $sp, $zero
        46 => x"AFC40008", -- sw $a0, 8(fp)
        47 => x"AFC5000C", -- sw $a1, 12(fp)
        48 => x"AFC60010", -- sw $a2, 16(fp)
        49 => x"0800003C", -- j 60
        50 => x"00000000", -- nop
        51 => x"8FC30008", -- lw $v1, 8(fp)
        52 => x"8FC2000C", -- lw $v0, 12(fp)
        53 => x"00000000", -- nop
        54 => x"304200FF", -- andi $v0, $v0, 00ff
        55 => x"A0620000", -- sb $v0, 0(v1)
        56 => x"8FC20008", -- lw $v0, 8(fp)
        57 => x"00000000", -- nop
        58 => x"24420001", -- addiu $v0, $v0, 1
        59 => x"AFC20008", -- sw $v0, 8(fp)
        60 => x"8FC20010", -- lw $v0, 16(fp)
        61 => x"00000000", -- nop
        62 => x"0002102B", -- sltu $v0, $zero, $v0
        63 => x"304300FF", -- andi $v1, $v0, 00ff
        64 => x"8FC20010", -- lw $v0, 16(fp)
        65 => x"00000000", -- nop
        66 => x"2442FFFF", -- addiu $v0, $v0, -1
        67 => x"AFC20010", -- sw $v0, 16(fp)
        68 => x"1460FFEE", -- bne $v1, $zero, -18
        69 => x"00000000", -- nop
        70 => x"03C0E821", -- addu $sp, $fp, $zero
        71 => x"8FBE0004", -- lw $fp, 4(sp)
        72 => x"27BD0008", -- addiu $sp, $sp, 8
        73 => x"03E00008", -- jr $ra
        74 => x"00000000", -- nop
        75 => x"27BDFFF0", -- addiu $sp, $sp, -16
        76 => x"AFBE000C", -- sw $fp, 12(sp)
        77 => x"03A0F021", -- addu $fp, $sp, $zero
        78 => x"AFC40010", -- sw $a0, 16(fp)
        79 => x"8FC20010", -- lw $v0, 16(fp)
        80 => x"00000000", -- nop
        81 => x"04410007", -- bgez $v0, 7
        82 => x"00000000", -- nop
        83 => x"8FC20010", -- lw $v0, 16(fp)
        84 => x"00000000", -- nop
        85 => x"00021023", -- subu $v0, $zero, $v0
        86 => x"AFC20000", -- sw $v0, 0(fp)
        87 => x"0800005C", -- j 92
        88 => x"00000000", -- nop
        89 => x"8FC20010", -- lw $v0, 16(fp)
        90 => x"00000000", -- nop
        91 => x"AFC20000", -- sw $v0, 0(fp)
        92 => x"8FC20000", -- lw $v0, 0(fp)
        93 => x"03C0E821", -- addu $sp, $fp, $zero
        94 => x"8FBE000C", -- lw $fp, 12(sp)
        95 => x"27BD0010", -- addiu $sp, $sp, 16
        96 => x"03E00008", -- jr $ra
        97 => x"00000000", -- nop
        98 => x"27BDFFD0", -- addiu $sp, $sp, -48
        99 => x"AFBF002C", -- sw $ra, 44(sp)
       100 => x"AFBE0028", -- sw $fp, 40(sp)
       101 => x"AFB10024", -- sw $s1, 36(sp)
       102 => x"AFB00020", -- sw $s0, 32(sp)
       103 => x"03A0F021", -- addu $fp, $sp, $zero
       104 => x"AFC40030", -- sw $a0, 48(fp)
       105 => x"AFC50034", -- sw $a1, 52(fp)
       106 => x"8F820850", -- lw $v0, 2128(gp)
       107 => x"8FC30034", -- lw $v1, 52(fp)
       108 => x"00000000", -- nop
       109 => x"0062102A", -- slt $v0, $v1, $v0
       110 => x"104000FB", -- beq $v0, $zero, 251
       111 => x"00000000", -- nop
       112 => x"8F83084C", -- lw $v1, 2124(gp)
       113 => x"8FC20030", -- lw $v0, 48(fp)
       114 => x"00000000", -- nop
       115 => x"14430006", -- bne $v0, $v1, 6
       116 => x"00000000", -- nop
       117 => x"8FC20034", -- lw $v0, 52(fp)
       118 => x"00000000", -- nop
       119 => x"AF820850", -- sw $v0, 2128(gp)
       120 => x"0800016A", -- j 362
       121 => x"00000000", -- nop
       122 => x"AFC0001C", -- sw $zero, 28(fp)
       123 => x"08000165", -- j 357
       124 => x"00000000", -- nop
       125 => x"AFC00018", -- sw $zero, 24(fp)
       126 => x"0800015C", -- j 348
       127 => x"00000000", -- nop
       128 => x"8FC20030", -- lw $v0, 48(fp)
       129 => x"00000000", -- nop
       130 => x"14400005", -- bne $v0, $zero, 5
       131 => x"00000000", -- nop
       132 => x"24020001", -- addiu $v0, $zero, 1
       133 => x"AFC20010", -- sw $v0, 16(fp)
       134 => x"080000F6", -- j 246
       135 => x"00000000", -- nop
       136 => x"8FC2001C", -- lw $v0, 28(fp)
       137 => x"8FC40018", -- lw $a0, 24(fp)
       138 => x"3C050000", -- lui $a1, 0000
       139 => x"00021040", -- sll $v0, $v0, 2
       140 => x"00021880", -- sll $v1, $v0, 4
       141 => x"00431021", -- addu $v0, $v0, $v1
       142 => x"00441021", -- addu $v0, $v0, $a0
       143 => x"00021880", -- sll $v1, $v0, 4
       144 => x"24A208B0", -- addiu $v0, $a1, 2224
       145 => x"00621021", -- addu $v0, $v1, $v0
       146 => x"8C420000", -- lw $v0, 0(v0)
       147 => x"00000000", -- nop
       148 => x"14400060", -- bne $v0, $zero, 96
       149 => x"00000000", -- nop
       150 => x"AFC00010", -- sw $zero, 16(fp)
       151 => x"8FC2001C", -- lw $v0, 28(fp)
       152 => x"00000000", -- nop
       153 => x"18400013", -- blez $v0, 19
       154 => x"00000000", -- nop
       155 => x"8FC2001C", -- lw $v0, 28(fp)
       156 => x"00000000", -- nop
       157 => x"2442FFFF", -- addiu $v0, $v0, -1
       158 => x"8FC40018", -- lw $a0, 24(fp)
       159 => x"3C050000", -- lui $a1, 0000
       160 => x"00021040", -- sll $v0, $v0, 2
       161 => x"00021880", -- sll $v1, $v0, 4
       162 => x"00431021", -- addu $v0, $v0, $v1
       163 => x"00441021", -- addu $v0, $v0, $a0
       164 => x"00021880", -- sll $v1, $v0, 4
       165 => x"24A208B0", -- addiu $v0, $a1, 2224
       166 => x"00621021", -- addu $v0, $v1, $v0
       167 => x"8C430000", -- lw $v1, 0(v0)
       168 => x"24020001", -- addiu $v0, $zero, 1
       169 => x"14620003", -- bne $v1, $v0, 3
       170 => x"00000000", -- nop
       171 => x"24020001", -- addiu $v0, $zero, 1
       172 => x"AFC20010", -- sw $v0, 16(fp)
       173 => x"8FC20018", -- lw $v0, 24(fp)
       174 => x"00000000", -- nop
       175 => x"18400014", -- blez $v0, 20
       176 => x"00000000", -- nop
       177 => x"8FC3001C", -- lw $v1, 28(fp)
       178 => x"8FC20018", -- lw $v0, 24(fp)
       179 => x"00000000", -- nop
       180 => x"2444FFFF", -- addiu $a0, $v0, -1
       181 => x"3C050000", -- lui $a1, 0000
       182 => x"00601021", -- addu $v0, $v1, $zero
       183 => x"00021040", -- sll $v0, $v0, 2
       184 => x"00021880", -- sll $v1, $v0, 4
       185 => x"00431021", -- addu $v0, $v0, $v1
       186 => x"00441021", -- addu $v0, $v0, $a0
       187 => x"00021880", -- sll $v1, $v0, 4
       188 => x"24A208B0", -- addiu $v0, $a1, 2224
       189 => x"00621021", -- addu $v0, $v1, $v0
       190 => x"8C430000", -- lw $v1, 0(v0)
       191 => x"24020001", -- addiu $v0, $zero, 1
       192 => x"14620003", -- bne $v1, $v0, 3
       193 => x"00000000", -- nop
       194 => x"24020001", -- addiu $v0, $zero, 1
       195 => x"AFC20010", -- sw $v0, 16(fp)
       196 => x"8FC2001C", -- lw $v0, 28(fp)
       197 => x"00000000", -- nop
       198 => x"28420004", -- slti $v0, $v0, 4
       199 => x"10400013", -- beq $v0, $zero, 19
       200 => x"00000000", -- nop
       201 => x"8FC2001C", -- lw $v0, 28(fp)
       202 => x"00000000", -- nop
       203 => x"24420001", -- addiu $v0, $v0, 1
       204 => x"8FC40018", -- lw $a0, 24(fp)
       205 => x"3C050000", -- lui $a1, 0000
       206 => x"00021040", -- sll $v0, $v0, 2
       207 => x"00021880", -- sll $v1, $v0, 4
       208 => x"00431021", -- addu $v0, $v0, $v1
       209 => x"00441021", -- addu $v0, $v0, $a0
       210 => x"00021880", -- sll $v1, $v0, 4
       211 => x"24A208B0", -- addiu $v0, $a1, 2224
       212 => x"00621021", -- addu $v0, $v1, $v0
       213 => x"8C430000", -- lw $v1, 0(v0)
       214 => x"24020001", -- addiu $v0, $zero, 1
       215 => x"14620003", -- bne $v1, $v0, 3
       216 => x"00000000", -- nop
       217 => x"24020001", -- addiu $v0, $zero, 1
       218 => x"AFC20010", -- sw $v0, 16(fp)
       219 => x"8FC20018", -- lw $v0, 24(fp)
       220 => x"00000000", -- nop
       221 => x"28420004", -- slti $v0, $v0, 4
       222 => x"10400017", -- beq $v0, $zero, 23
       223 => x"00000000", -- nop
       224 => x"8FC3001C", -- lw $v1, 28(fp)
       225 => x"8FC20018", -- lw $v0, 24(fp)
       226 => x"00000000", -- nop
       227 => x"24440001", -- addiu $a0, $v0, 1
       228 => x"3C050000", -- lui $a1, 0000
       229 => x"00601021", -- addu $v0, $v1, $zero
       230 => x"00021040", -- sll $v0, $v0, 2
       231 => x"00021880", -- sll $v1, $v0, 4
       232 => x"00431021", -- addu $v0, $v0, $v1
       233 => x"00441021", -- addu $v0, $v0, $a0
       234 => x"00021880", -- sll $v1, $v0, 4
       235 => x"24A208B0", -- addiu $v0, $a1, 2224
       236 => x"00621021", -- addu $v0, $v1, $v0
       237 => x"8C430000", -- lw $v1, 0(v0)
       238 => x"24020001", -- addiu $v0, $zero, 1
       239 => x"14620006", -- bne $v1, $v0, 6
       240 => x"00000000", -- nop
       241 => x"24020001", -- addiu $v0, $zero, 1
       242 => x"AFC20010", -- sw $v0, 16(fp)
       243 => x"080000F6", -- j 246
       244 => x"00000000", -- nop
       245 => x"AFC00010", -- sw $zero, 16(fp)
       246 => x"8FC20010", -- lw $v0, 16(fp)
       247 => x"00000000", -- nop
       248 => x"1040005F", -- beq $v0, $zero, 95
       249 => x"00000000", -- nop
       250 => x"8FC2001C", -- lw $v0, 28(fp)
       251 => x"8FC40018", -- lw $a0, 24(fp)
       252 => x"3C050000", -- lui $a1, 0000
       253 => x"00021040", -- sll $v0, $v0, 2
       254 => x"00021880", -- sll $v1, $v0, 4
       255 => x"00431021", -- addu $v0, $v0, $v1
       256 => x"00441021", -- addu $v0, $v0, $a0
       257 => x"00021880", -- sll $v1, $v0, 4
       258 => x"24A208B0", -- addiu $v0, $a1, 2224
       259 => x"00621821", -- addu $v1, $v1, $v0
       260 => x"24020001", -- addiu $v0, $zero, 1
       261 => x"AC620000", -- sw $v0, 0(v1)
       262 => x"AFC00014", -- sw $zero, 20(fp)
       263 => x"08000147", -- j 327
       264 => x"00000000", -- nop
       265 => x"8FC20014", -- lw $v0, 20(fp)
       266 => x"3C030000", -- lui $v1, 0000
       267 => x"00022080", -- sll $a0, $v0, 4
       268 => x"24620A40", -- addiu $v0, $v1, 2624
       269 => x"00821021", -- addu $v0, $a0, $v0
       270 => x"8C420000", -- lw $v0, 0(v0)
       271 => x"00000000", -- nop
       272 => x"14400032", -- bne $v0, $zero, 50
       273 => x"00000000", -- nop
       274 => x"8FC20014", -- lw $v0, 20(fp)
       275 => x"3C030000", -- lui $v1, 0000
       276 => x"00022080", -- sll $a0, $v0, 4
       277 => x"24620A40", -- addiu $v0, $v1, 2624
       278 => x"00821821", -- addu $v1, $a0, $v0
       279 => x"24020001", -- addiu $v0, $zero, 1
       280 => x"AC620000", -- sw $v0, 0(v1)
       281 => x"8FC20030", -- lw $v0, 48(fp)
       282 => x"00000000", -- nop
       283 => x"24500001", -- addiu $s0, $v0, 1
       284 => x"8FC20014", -- lw $v0, 20(fp)
       285 => x"3C030000", -- lui $v1, 0000
       286 => x"00022080", -- sll $a0, $v0, 4
       287 => x"24620854", -- addiu $v0, $v1, 2132
       288 => x"00821021", -- addu $v0, $a0, $v0
       289 => x"8C430000", -- lw $v1, 0(v0)
       290 => x"8FC2001C", -- lw $v0, 28(fp)
       291 => x"00000000", -- nop
       292 => x"00621023", -- subu $v0, $v1, $v0
       293 => x"00402021", -- addu $a0, $v0, $zero
       294 => x"0C00004B", -- jal 75
       295 => x"00000000", -- nop
       296 => x"00401821", -- addu $v1, $v0, $zero
       297 => x"8FC20034", -- lw $v0, 52(fp)
       298 => x"00000000", -- nop
       299 => x"00628821", -- addu $s1, $v1, $v0
       300 => x"8FC20014", -- lw $v0, 20(fp)
       301 => x"3C030000", -- lui $v1, 0000
       302 => x"00022080", -- sll $a0, $v0, 4
       303 => x"24620888", -- addiu $v0, $v1, 2184
       304 => x"00821021", -- addu $v0, $a0, $v0
       305 => x"8C430000", -- lw $v1, 0(v0)
       306 => x"8FC20018", -- lw $v0, 24(fp)
       307 => x"00000000", -- nop
       308 => x"00621023", -- subu $v0, $v1, $v0
       309 => x"00402021", -- addu $a0, $v0, $zero
       310 => x"0C00004B", -- jal 75
       311 => x"00000000", -- nop
       312 => x"02221021", -- addu $v0, $s1, $v0
       313 => x"02002021", -- addu $a0, $s0, $zero
       314 => x"00402821", -- addu $a1, $v0, $zero
       315 => x"0C000062", -- jal 98
       316 => x"00000000", -- nop
       317 => x"8FC20014", -- lw $v0, 20(fp)
       318 => x"3C030000", -- lui $v1, 0000
       319 => x"00022080", -- sll $a0, $v0, 4
       320 => x"24620A40", -- addiu $v0, $v1, 2624
       321 => x"00821021", -- addu $v0, $a0, $v0
       322 => x"AC400000", -- sw $zero, 0(v0)
       323 => x"8FC20014", -- lw $v0, 20(fp)
       324 => x"00000000", -- nop
       325 => x"24420001", -- addiu $v0, $v0, 1
       326 => x"AFC20014", -- sw $v0, 20(fp)
       327 => x"8F82084C", -- lw $v0, 2124(gp)
       328 => x"8FC30014", -- lw $v1, 20(fp)
       329 => x"00000000", -- nop
       330 => x"0062102A", -- slt $v0, $v1, $v0
       331 => x"1440FFBD", -- bne $v0, $zero, -67
       332 => x"00000000", -- nop
       333 => x"8FC2001C", -- lw $v0, 28(fp)
       334 => x"8FC40018", -- lw $a0, 24(fp)
       335 => x"3C050000", -- lui $a1, 0000
       336 => x"00021040", -- sll $v0, $v0, 2
       337 => x"00021880", -- sll $v1, $v0, 4
       338 => x"00431021", -- addu $v0, $v0, $v1
       339 => x"00441021", -- addu $v0, $v0, $a0
       340 => x"00021880", -- sll $v1, $v0, 4
       341 => x"24A208B0", -- addiu $v0, $a1, 2224
       342 => x"00621021", -- addu $v0, $v1, $v0
       343 => x"AC400000", -- sw $zero, 0(v0)
       344 => x"8FC20018", -- lw $v0, 24(fp)
       345 => x"00000000", -- nop
       346 => x"24420001", -- addiu $v0, $v0, 1
       347 => x"AFC20018", -- sw $v0, 24(fp)
       348 => x"8FC20018", -- lw $v0, 24(fp)
       349 => x"00000000", -- nop
       350 => x"28420005", -- slti $v0, $v0, 5
       351 => x"1440FF20", -- bne $v0, $zero, -224
       352 => x"00000000", -- nop
       353 => x"8FC2001C", -- lw $v0, 28(fp)
       354 => x"00000000", -- nop
       355 => x"24420001", -- addiu $v0, $v0, 1
       356 => x"AFC2001C", -- sw $v0, 28(fp)
       357 => x"8FC2001C", -- lw $v0, 28(fp)
       358 => x"00000000", -- nop
       359 => x"28420005", -- slti $v0, $v0, 5
       360 => x"1440FF14", -- bne $v0, $zero, -236
       361 => x"00000000", -- nop
       362 => x"03C0E821", -- addu $sp, $fp, $zero
       363 => x"8FBF002C", -- lw $ra, 44(sp)
       364 => x"8FBE0028", -- lw $fp, 40(sp)
       365 => x"8FB10024", -- lw $s1, 36(sp)
       366 => x"8FB00020", -- lw $s0, 32(sp)
       367 => x"27BD0030", -- addiu $sp, $sp, 48
       368 => x"03E00008", -- jr $ra
       369 => x"00000000", -- nop
       370 => x"27BDFFE0", -- addiu $sp, $sp, -32
       371 => x"AFBF001C", -- sw $ra, 28(sp)
       372 => x"AFBE0018", -- sw $fp, 24(sp)
       373 => x"03A0F021", -- addu $fp, $sp, $zero
       374 => x"AFC40020", -- sw $a0, 32(fp)
       375 => x"AF80084C", -- sw $zero, 2124(gp)
       376 => x"AFC00014", -- sw $zero, 20(fp)
       377 => x"080001AE", -- j 430
       378 => x"00000000", -- nop
       379 => x"AFC00010", -- sw $zero, 16(fp)
       380 => x"080001A5", -- j 421
       381 => x"00000000", -- nop
       382 => x"8FC30014", -- lw $v1, 20(fp)
       383 => x"00000000", -- nop
       384 => x"00601021", -- addu $v0, $v1, $zero
       385 => x"00021080", -- sll $v0, $v0, 4
       386 => x"00431821", -- addu $v1, $v0, $v1
       387 => x"8FC20020", -- lw $v0, 32(fp)
       388 => x"00000000", -- nop
       389 => x"00431821", -- addu $v1, $v0, $v1
       390 => x"8FC20010", -- lw $v0, 16(fp)
       391 => x"00000000", -- nop
       392 => x"00621021", -- addu $v0, $v1, $v0
       393 => x"80430000", -- lb $v1, 0(v0)
       394 => x"2402002A", -- addiu $v0, $zero, 42
       395 => x"14620015", -- bne $v1, $v0, 21
       396 => x"00000000", -- nop
       397 => x"8F82084C", -- lw $v0, 2124(gp)
       398 => x"3C030000", -- lui $v1, 0000
       399 => x"00022080", -- sll $a0, $v0, 4
       400 => x"24620854", -- addiu $v0, $v1, 2132
       401 => x"00821821", -- addu $v1, $a0, $v0
       402 => x"8FC20014", -- lw $v0, 20(fp)
       403 => x"00000000", -- nop
       404 => x"AC620000", -- sw $v0, 0(v1)
       405 => x"8F82084C", -- lw $v0, 2124(gp)
       406 => x"3C030000", -- lui $v1, 0000
       407 => x"00022080", -- sll $a0, $v0, 4
       408 => x"24620888", -- addiu $v0, $v1, 2184
       409 => x"00821821", -- addu $v1, $a0, $v0
       410 => x"8FC20010", -- lw $v0, 16(fp)
       411 => x"00000000", -- nop
       412 => x"AC620000", -- sw $v0, 0(v1)
       413 => x"8F82084C", -- lw $v0, 2124(gp)
       414 => x"00000000", -- nop
       415 => x"24420001", -- addiu $v0, $v0, 1
       416 => x"AF82084C", -- sw $v0, 2124(gp)
       417 => x"8FC20010", -- lw $v0, 16(fp)
       418 => x"00000000", -- nop
       419 => x"24420001", -- addiu $v0, $v0, 1
       420 => x"AFC20010", -- sw $v0, 16(fp)
       421 => x"8FC20010", -- lw $v0, 16(fp)
       422 => x"00000000", -- nop
       423 => x"28420005", -- slti $v0, $v0, 5
       424 => x"1440FFD5", -- bne $v0, $zero, -43
       425 => x"00000000", -- nop
       426 => x"8FC20014", -- lw $v0, 20(fp)
       427 => x"00000000", -- nop
       428 => x"24420001", -- addiu $v0, $v0, 1
       429 => x"AFC20014", -- sw $v0, 20(fp)
       430 => x"8FC20014", -- lw $v0, 20(fp)
       431 => x"00000000", -- nop
       432 => x"28420005", -- slti $v0, $v0, 5
       433 => x"1440FFC9", -- bne $v0, $zero, -55
       434 => x"00000000", -- nop
       435 => x"3C020000", -- lui $v0, 0000
       436 => x"244408B0", -- addiu $a0, $v0, 2224
       437 => x"00002821", -- addu $a1, $zero, $zero
       438 => x"24060190", -- addiu $a2, $zero, 400
       439 => x"0C00002B", -- jal 43
       440 => x"00000000", -- nop
       441 => x"3C020000", -- lui $v0, 0000
       442 => x"24440A40", -- addiu $a0, $v0, 2624
       443 => x"00002821", -- addu $a1, $zero, $zero
       444 => x"24060028", -- addiu $a2, $zero, 40
       445 => x"0C00002B", -- jal 43
       446 => x"00000000", -- nop
       447 => x"3C02000F", -- lui $v0, 000f
       448 => x"34424240", -- ori $v0, $v0, 4240
       449 => x"AF820850", -- sw $v0, 2128(gp)
       450 => x"00002021", -- addu $a0, $zero, $zero
       451 => x"00002821", -- addu $a1, $zero, $zero
       452 => x"0C000062", -- jal 98
       453 => x"00000000", -- nop
       454 => x"8F820850", -- lw $v0, 2128(gp)
       455 => x"03C0E821", -- addu $sp, $fp, $zero
       456 => x"8FBF001C", -- lw $ra, 28(sp)
       457 => x"8FBE0018", -- lw $fp, 24(sp)
       458 => x"27BD0020", -- addiu $sp, $sp, 32
       459 => x"03E00008", -- jr $ra
       460 => x"00000000", -- nop
       461 => x"27BDFFD8", -- addiu $sp, $sp, -40
       462 => x"AFBF0024", -- sw $ra, 36(sp)
       463 => x"AFBE0020", -- sw $fp, 32(sp)
       464 => x"AFB0001C", -- sw $s0, 28(sp)
       465 => x"03A0F021", -- addu $fp, $sp, $zero
       466 => x"AFC00010", -- sw $zero, 16(fp)
       467 => x"080001ED", -- j 493
       468 => x"00000000", -- nop
       469 => x"8FD00010", -- lw $s0, 16(fp)
       470 => x"3C020000", -- lui $v0, 0000
       471 => x"24450800", -- addiu $a1, $v0, 2048
       472 => x"8FC40010", -- lw $a0, 16(fp)
       473 => x"00000000", -- nop
       474 => x"00801021", -- addu $v0, $a0, $zero
       475 => x"000218C0", -- sll $v1, $v0, 6
       476 => x"00031080", -- sll $v0, $v1, 4
       477 => x"00431023", -- subu $v0, $v0, $v1
       478 => x"00441021", -- addu $v0, $v0, $a0
       479 => x"00A21021", -- addu $v0, $a1, $v0
       480 => x"00402021", -- addu $a0, $v0, $zero
       481 => x"0C000172", -- jal 370
       482 => x"00000000", -- nop
       483 => x"00402021", -- addu $a0, $v0, $zero
       484 => x"3C020000", -- lui $v0, 0000
       485 => x"00101880", -- sll $v1, $s0, 4
       486 => x"2442087C", -- addiu $v0, $v0, 2172
       487 => x"00621021", -- addu $v0, $v1, $v0
       488 => x"AC440000", -- sw $a0, 0(v0)
       489 => x"8FC20010", -- lw $v0, 16(fp)
       490 => x"00000000", -- nop
       491 => x"24420001", -- addiu $v0, $v0, 1
       492 => x"AFC20010", -- sw $v0, 16(fp)
       493 => x"8FC20010", -- lw $v0, 16(fp)
       494 => x"00000000", -- nop
       495 => x"28420003", -- slti $v0, $v0, 3
       496 => x"1440FFE4", -- bne $v0, $zero, -28
       497 => x"00000000", -- nop
       498 => x"00001021", -- addu $v0, $zero, $zero
       499 => x"03C0E821", -- addu $sp, $fp, $zero
       500 => x"8FBF0024", -- lw $ra, 36(sp)
       501 => x"8FBE0020", -- lw $fp, 32(sp)
       502 => x"8FB0001C", -- lw $s0, 28(sp)
       503 => x"27BD0028", -- addiu $sp, $sp, 40
       504 => x"03E00008", -- jr $ra
       505 => x"00000000", -- nop
       506 => x"00000000", -- nop
       507 => x"00000000", -- nop
       508 => x"00000000", -- nop
       509 => x"00000000", -- nop
       510 => x"00000000", -- nop
       511 => x"00000000"  -- nop
    );

BEGIN

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF R='1' THEN
                DATA_OUT <= TMP_RAM(CONV_INTEGER(UNSIGNED(RADDR(ADDR-1 DOWNTO 2))));
            ELSE
                DATA_OUT <= (DATA_OUT'RANGE => 'Z');
            END IF;
        END IF;
    END IF;
    END PROCESS;

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF W='1' THEN
                TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2)))) <= DATA_IN;
            END IF;
        END IF;
    END IF;
    END PROCESS;

END BEHAV_CODE;

ARCHITECTURE BEHAV_DATA OF SRAM IS

    TYPE RAM_TYPE IS ARRAY (0 TO DEPTH-1) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL IBYTE0:     STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL IBYTE1:     STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL IBYTE2:     STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL IBYTE3:     STD_LOGIC_VECTOR(7 DOWNTO 0);

    SIGNAL OBYTE:      STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL OHALF:      STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SBYTE:      STD_LOGIC_VECTOR(23 DOWNTO 0);
    SIGNAL SHALF:      STD_LOGIC_VECTOR(15 DOWNTO 0);

    SIGNAL RWORD:      STD_LOGIC_VECTOR(31 DOWNTO 0):= x"00000000";

    SIGNAL RADDR2:     STD_LOGIC_VECTOR(1 DOWNTO 0):= "00";
    SIGNAL MODE2:      STD_LOGIC_VECTOR(2 DOWNTO 0):= "000";
    SIGNAL ISSIGNED2:  STD_LOGIC:= '0';

    SIGNAL W0:         STD_LOGIC;
    SIGNAL W1:         STD_LOGIC;
    SIGNAL W2:         STD_LOGIC;
    SIGNAL W3:         STD_LOGIC;

    SIGNAL TMP_RAM: RAM_TYPE := (

         0 => x"2E2E2E2E",
         1 => x"2E2E2E2A",
         2 => x"2A2E2E2E",
         3 => x"2E2E2E2E",
         4 => x"2E2E2A2E",
         5 => x"2E2E2E2E",
         6 => x"2E2E2E2E",
         7 => x"2E2E2E2E",
         8 => x"2E2E2E2E",
         9 => x"2A2A2E2E",
        10 => x"2E2A2E2E",
        11 => x"2E2A2A2E",
        12 => x"2E2E2A2E",
        13 => x"2E2E2A2E",
        14 => x"2E2E2E2E",
        15 => x"2E2E2E2E",
        16 => x"2E2E2E2E",
        17 => x"2E2E2A2E",
        18 => x"2E2E2A00",
        19 => x"55555555",
        20 => x"55555555",
        21 => x"55555555",
        22 => x"55555555",
        23 => x"55555555",
        24 => x"55555555",
        25 => x"55555555",
        26 => x"55555555",
        27 => x"55555555",
        28 => x"55555555",
        29 => x"55555555",
        30 => x"55555555",
        31 => x"55555555",
        32 => x"55555555",
        33 => x"55555555",
        34 => x"55555555",
        35 => x"55555555",
        36 => x"55555555",
        37 => x"55555555",
        38 => x"55555555",
        39 => x"55555555",
        40 => x"55555555",
        41 => x"55555555",
        42 => x"55555555",
        43 => x"55555555",
        44 => x"55555555",
        45 => x"55555555",
        46 => x"55555555",
        47 => x"55555555",
        48 => x"55555555",
        49 => x"55555555",
        50 => x"55555555",
        51 => x"55555555",
        52 => x"55555555",
        53 => x"55555555",
        54 => x"55555555",
        55 => x"55555555",
        56 => x"55555555",
        57 => x"55555555",
        58 => x"55555555",
        59 => x"55555555",
        60 => x"55555555",
        61 => x"55555555",
        62 => x"55555555",
        63 => x"55555555",
        64 => x"55555555",
        65 => x"55555555",
        66 => x"55555555",
        67 => x"55555555",
        68 => x"55555555",
        69 => x"55555555",
        70 => x"55555555",
        71 => x"55555555",
        72 => x"55555555",
        73 => x"55555555",
        74 => x"55555555",
        75 => x"55555555",
        76 => x"55555555",
        77 => x"55555555",
        78 => x"55555555",
        79 => x"55555555",
        80 => x"55555555",
        81 => x"55555555",
        82 => x"55555555",
        83 => x"55555555",
        84 => x"55555555",
        85 => x"55555555",
        86 => x"55555555",
        87 => x"55555555",
        88 => x"55555555",
        89 => x"55555555",
        90 => x"55555555",
        91 => x"55555555",
        92 => x"55555555",
        93 => x"55555555",
        94 => x"55555555",
        95 => x"55555555",
        96 => x"55555555",
        97 => x"55555555",
        98 => x"55555555",
        99 => x"55555555",
       100 => x"55555555",
       101 => x"55555555",
       102 => x"55555555",
       103 => x"55555555",
       104 => x"55555555",
       105 => x"55555555",
       106 => x"55555555",
       107 => x"55555555",
       108 => x"55555555",
       109 => x"55555555",
       110 => x"55555555",
       111 => x"55555555",
       112 => x"55555555",
       113 => x"55555555",
       114 => x"55555555",
       115 => x"55555555",
       116 => x"55555555",
       117 => x"55555555",
       118 => x"55555555",
       119 => x"55555555",
       120 => x"55555555",
       121 => x"55555555",
       122 => x"55555555",
       123 => x"55555555",
       124 => x"55555555",
       125 => x"55555555",
       126 => x"55555555",
       127 => x"55555555",
       128 => x"55555555",
       129 => x"55555555",
       130 => x"55555555",
       131 => x"55555555",
       132 => x"55555555",
       133 => x"55555555",
       134 => x"55555555",
       135 => x"55555555",
       136 => x"55555555",
       137 => x"55555555",
       138 => x"55555555",
       139 => x"55555555",
       140 => x"55555555",
       141 => x"55555555",
       142 => x"55555555",
       143 => x"55555555",
       144 => x"55555555",
       145 => x"55555555",
       146 => x"55555555",
       147 => x"55555555",
       148 => x"55555555",
       149 => x"55555555",
       150 => x"55555555",
       151 => x"55555555",
       152 => x"55555555",
       153 => x"55555555",
       154 => x"55555555",
       155 => x"55555555",
       156 => x"55555555",
       157 => x"55555555",
       158 => x"55555555",
       159 => x"55555555",
       160 => x"55555555",
       161 => x"55555555",
       162 => x"55555555",
       163 => x"55555555",
       164 => x"55555555",
       165 => x"55555555",
       166 => x"55555555",
       167 => x"55555555",
       168 => x"55555555",
       169 => x"55555555",
       170 => x"55555555",
       171 => x"55555555",
       172 => x"55555555",
       173 => x"55555555",
       174 => x"55555555",
       175 => x"55555555",
       176 => x"55555555",
       177 => x"55555555",
       178 => x"55555555",
       179 => x"55555555",
       180 => x"55555555",
       181 => x"55555555",
       182 => x"55555555",
       183 => x"55555555",
       184 => x"55555555",
       185 => x"55555555",
       186 => x"55555555",
       187 => x"55555555",
       188 => x"55555555",
       189 => x"55555555",
       190 => x"55555555",
       191 => x"55555555",
       192 => x"55555555",
       193 => x"55555555",
       194 => x"55555555",
       195 => x"55555555",
       196 => x"55555555",
       197 => x"55555555",
       198 => x"55555555",
       199 => x"55555555",
       200 => x"55555555",
       201 => x"55555555",
       202 => x"55555555",
       203 => x"55555555",
       204 => x"55555555",
       205 => x"55555555",
       206 => x"55555555",
       207 => x"55555555",
       208 => x"55555555",
       209 => x"55555555",
       210 => x"55555555",
       211 => x"55555555",
       212 => x"55555555",
       213 => x"55555555",
       214 => x"55555555",
       215 => x"55555555",
       216 => x"55555555",
       217 => x"55555555",
       218 => x"55555555",
       219 => x"55555555",
       220 => x"55555555",
       221 => x"55555555",
       222 => x"55555555",
       223 => x"55555555",
       224 => x"55555555",
       225 => x"55555555",
       226 => x"55555555",
       227 => x"55555555",
       228 => x"55555555",
       229 => x"55555555",
       230 => x"55555555",
       231 => x"55555555",
       232 => x"55555555",
       233 => x"55555555",
       234 => x"55555555",
       235 => x"55555555",
       236 => x"55555555",
       237 => x"55555555",
       238 => x"55555555",
       239 => x"55555555",
       240 => x"55555555",
       241 => x"55555555",
       242 => x"55555555",
       243 => x"55555555",
       244 => x"55555555",
       245 => x"55555555",
       246 => x"55555555",
       247 => x"55555555",
       248 => x"55555555",
       249 => x"55555555",
       250 => x"55555555",
       251 => x"55555555",
       252 => x"55555555",
       253 => x"55555555",
       254 => x"55555555",
       255 => x"55555555",
       256 => x"55555555",
       257 => x"55555555",
       258 => x"55555555",
       259 => x"55555555",
       260 => x"55555555",
       261 => x"55555555",
       262 => x"55555555",
       263 => x"55555555",
       264 => x"55555555",
       265 => x"55555555",
       266 => x"55555555",
       267 => x"55555555",
       268 => x"55555555",
       269 => x"55555555",
       270 => x"55555555",
       271 => x"55555555",
       272 => x"55555555",
       273 => x"55555555",
       274 => x"55555555",
       275 => x"55555555",
       276 => x"55555555",
       277 => x"55555555",
       278 => x"55555555",
       279 => x"55555555",
       280 => x"55555555",
       281 => x"55555555",
       282 => x"55555555",
       283 => x"55555555",
       284 => x"55555555",
       285 => x"55555555",
       286 => x"55555555",
       287 => x"55555555",
       288 => x"55555555",
       289 => x"55555555",
       290 => x"55555555",
       291 => x"55555555",
       292 => x"55555555",
       293 => x"55555555",
       294 => x"55555555",
       295 => x"55555555",
       296 => x"55555555",
       297 => x"55555555",
       298 => x"55555555",
       299 => x"55555555",
       300 => x"55555555",
       301 => x"55555555",
       302 => x"55555555",
       303 => x"55555555",
       304 => x"55555555",
       305 => x"55555555",
       306 => x"55555555",
       307 => x"55555555",
       308 => x"55555555",
       309 => x"55555555",
       310 => x"55555555",
       311 => x"55555555",
       312 => x"55555555",
       313 => x"55555555",
       314 => x"55555555",
       315 => x"55555555",
       316 => x"55555555",
       317 => x"55555555",
       318 => x"55555555",
       319 => x"55555555",
       320 => x"55555555",
       321 => x"55555555",
       322 => x"55555555",
       323 => x"55555555",
       324 => x"55555555",
       325 => x"55555555",
       326 => x"55555555",
       327 => x"55555555",
       328 => x"55555555",
       329 => x"55555555",
       330 => x"55555555",
       331 => x"55555555",
       332 => x"55555555",
       333 => x"55555555",
       334 => x"55555555",
       335 => x"55555555",
       336 => x"55555555",
       337 => x"55555555",
       338 => x"55555555",
       339 => x"55555555",
       340 => x"55555555",
       341 => x"55555555",
       342 => x"55555555",
       343 => x"55555555",
       344 => x"55555555",
       345 => x"55555555",
       346 => x"55555555",
       347 => x"55555555",
       348 => x"55555555",
       349 => x"55555555",
       350 => x"55555555",
       351 => x"55555555",
       352 => x"55555555",
       353 => x"55555555",
       354 => x"55555555",
       355 => x"55555555",
       356 => x"55555555",
       357 => x"55555555",
       358 => x"55555555",
       359 => x"55555555",
       360 => x"55555555",
       361 => x"55555555",
       362 => x"55555555",
       363 => x"55555555",
       364 => x"55555555",
       365 => x"55555555",
       366 => x"55555555",
       367 => x"55555555",
       368 => x"55555555",
       369 => x"55555555",
       370 => x"55555555",
       371 => x"55555555",
       372 => x"55555555",
       373 => x"55555555",
       374 => x"55555555",
       375 => x"55555555",
       376 => x"55555555",
       377 => x"55555555",
       378 => x"55555555",
       379 => x"55555555",
       380 => x"55555555",
       381 => x"55555555",
       382 => x"55555555",
       383 => x"55555555",
       384 => x"55555555",
       385 => x"55555555",
       386 => x"55555555",
       387 => x"55555555",
       388 => x"55555555",
       389 => x"55555555",
       390 => x"55555555",
       391 => x"55555555",
       392 => x"55555555",
       393 => x"55555555",
       394 => x"55555555",
       395 => x"55555555",
       396 => x"55555555",
       397 => x"55555555",
       398 => x"55555555",
       399 => x"55555555",
       400 => x"55555555",
       401 => x"55555555",
       402 => x"55555555",
       403 => x"55555555",
       404 => x"55555555",
       405 => x"55555555",
       406 => x"55555555",
       407 => x"55555555",
       408 => x"55555555",
       409 => x"55555555",
       410 => x"55555555",
       411 => x"55555555",
       412 => x"55555555",
       413 => x"55555555",
       414 => x"55555555",
       415 => x"55555555",
       416 => x"55555555",
       417 => x"55555555",
       418 => x"55555555",
       419 => x"55555555",
       420 => x"55555555",
       421 => x"55555555",
       422 => x"55555555",
       423 => x"55555555",
       424 => x"55555555",
       425 => x"55555555",
       426 => x"55555555",
       427 => x"55555555",
       428 => x"55555555",
       429 => x"55555555",
       430 => x"55555555",
       431 => x"55555555",
       432 => x"55555555",
       433 => x"55555555",
       434 => x"55555555",
       435 => x"55555555",
       436 => x"55555555",
       437 => x"55555555",
       438 => x"55555555",
       439 => x"55555555",
       440 => x"55555555",
       441 => x"55555555",
       442 => x"55555555",
       443 => x"55555555",
       444 => x"55555555",
       445 => x"55555555",
       446 => x"55555555",
       447 => x"55555555",
       448 => x"55555555",
       449 => x"55555555",
       450 => x"55555555",
       451 => x"55555555",
       452 => x"55555555",
       453 => x"55555555",
       454 => x"55555555",
       455 => x"55555555",
       456 => x"55555555",
       457 => x"55555555",
       458 => x"55555555",
       459 => x"55555555",
       460 => x"55555555",
       461 => x"55555555",
       462 => x"55555555",
       463 => x"55555555",
       464 => x"55555555",
       465 => x"55555555",
       466 => x"55555555",
       467 => x"55555555",
       468 => x"55555555",
       469 => x"55555555",
       470 => x"55555555",
       471 => x"55555555",
       472 => x"55555555",
       473 => x"55555555",
       474 => x"55555555",
       475 => x"55555555",
       476 => x"55555555",
       477 => x"55555555",
       478 => x"55555555",
       479 => x"55555555",
       480 => x"55555555",
       481 => x"55555555",
       482 => x"55555555",
       483 => x"55555555",
       484 => x"55555555",
       485 => x"55555555",
       486 => x"55555555",
       487 => x"55555555",
       488 => x"55555555",
       489 => x"55555555",
       490 => x"55555555",
       491 => x"55555555",
       492 => x"55555555",
       493 => x"55555555",
       494 => x"55555555",
       495 => x"55555555",
       496 => x"55555555",
       497 => x"55555555",
       498 => x"55555555",
       499 => x"55555555",
       500 => x"55555555",
       501 => x"55555555",
       502 => x"55555555",
       503 => x"55555555",
       504 => x"55555555",
       505 => x"55555555",
       506 => x"55555555",
       507 => x"55555555",
       508 => x"55555555",
       509 => x"55555555",
       510 => x"55555555",
       511 => x"55555555"
    );

BEGIN
    -- READ LOGIC
    OBYTE    <=      RWORD(31 DOWNTO 24) WHEN RADDR2(1 DOWNTO 0) = "00"
                ELSE RWORD(23 DOWNTO 16) WHEN RADDR2(1 DOWNTO 0) = "01"
                ELSE RWORD(15 DOWNTO  8) WHEN RADDR2(1 DOWNTO 0) = "10"
                ELSE RWORD( 7 DOWNTO  0);

    OHALF    <=      RWORD(31 DOWNTO 16) WHEN RADDR2(1 DOWNTO 0) = "00"
                ELSE RWORD(15 DOWNTO  0); -- THIS IS CASE "11", WE DON'T HANDLE THE OTHER CASES


    SBYTE    <=      x"FFFFFF" WHEN (OBYTE(7)  AND ISSIGNED2) = '1' ELSE x"000000";
    SHALF    <=      x"FFFF"   WHEN (OHALF(15) AND ISSIGNED2) = '1' ELSE x"0000";


    DATA_OUT <=      SBYTE & OBYTE WHEN MODE2(2) = '1'
                ELSE SHALF & OHALF WHEN MODE2(1) = '1'
                ELSE RWORD WHEN MODE2(0) = '1';

    -- WRITE LOGIC

    IBYTE0 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN(15 DOWNTO 8) WHEN MODE(1)='1' ELSE DATA_IN(31 DOWNTO  24);
    IBYTE1 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN( 7 DOWNTO 0) WHEN MODE(1)='1' ELSE DATA_IN(23 DOWNTO  16);
    IBYTE2 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN(15 DOWNTO 8) WHEN MODE(1)='1' ELSE DATA_IN(15 DOWNTO   8);
    IBYTE3 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN( 7 DOWNTO 0) WHEN MODE(1)='1' ELSE DATA_IN( 7 DOWNTO   0);

    W0 <= (   (MODE(2) AND NOT(WADDR(1) OR   WADDR(0)))  --B: "00"
           OR (MODE(1) AND NOT(WADDR(1)))                --H: "0x"
           OR  MODE(0)) AND W;                           --W: "Xx"
    W1 <= (   (MODE(2) AND NOT(WADDR(1)) AND WADDR(0))   --B: "01"
           OR (MODE(1) AND NOT(WADDR(1)))                --H: "0x"
           OR  MODE(0)) AND W;                           --W: "Xx"
    W2 <= (   (MODE(2) AND NOT(WADDR(0)) AND WADDR(1))   --B: "10"
           OR (MODE(1) AND     WADDR(1))                 --H: "1x"
           OR  MODE(0)) AND W;                           --W: "Xx"
    W3 <= (   (MODE(2) AND     WADDR(1) AND  WADDR(0))   --B: "11"
           OR (MODE(1) AND     WADDR(1))                 --H: "1x"
           OR  MODE(0)) AND W;                           --W: "Xx"

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        MODE2     <= MODE;
        ISSIGNED2 <= ISSIGNED;
        RADDR2 <= RADDR(1 DOWNTO 0);
    END IF;
    END PROCESS;

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF R='1' THEN
                RWORD <= TMP_RAM(CONV_INTEGER(UNSIGNED(RADDR(ADDR-1 DOWNTO 2))));
            ELSE
                RWORD <= (DATA_OUT'RANGE => 'Z');
            END IF;
        END IF;
    END IF;
    END PROCESS;

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF W='1' THEN
                IF W0 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(31 DOWNTO 24) <= IBYTE0;
                END IF;
                IF W1 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(23 DOWNTO 16) <= IBYTE1;
                END IF;
                IF W2 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(15 DOWNTO  8) <= IBYTE2;
                END IF;
                IF W3 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(7  DOWNTO  0) <= IBYTE3;
                END IF;
            END IF;
        END IF;
    END IF;
    END PROCESS;

END BEHAV_DATA;
