----------------------------------------------------------
--
-- 32 bits pipelined RISC processor
-- Copyright (c) 2010 Victor Munoz. All rights reserved.
-- derechos reservados, prohibida su reproduccion
--
-- Author: Victor Munoz
-- Contact: vmunoz@ingenieria-inversa.cl
--
----------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

----------------------------------------------------------

ENTITY SRAM IS
    GENERIC(
        ADDR:     INTEGER:= (9+2);
        DEPTH:    INTEGER:= 512
    );
    PORT(
        CLK:      IN  STD_LOGIC;
        ENABLE:   IN  STD_LOGIC;
        R:        IN  STD_LOGIC;
        W:        IN  STD_LOGIC;
        RADDR:    IN  STD_LOGIC_VECTOR(ADDR-1 DOWNTO 0);
        WADDR:    IN  STD_LOGIC_VECTOR(ADDR-1 DOWNTO 0);
        DATA_IN:  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
        MODE:     IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
        ISSIGNED: IN  STD_LOGIC;
        DATA_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0):= "00000000000000000000000000000000"
    );
END SRAM;

--------------------------------------------------------------

ARCHITECTURE BEHAV_CODE OF SRAM IS

    TYPE RAM_TYPE IS ARRAY (0 TO DEPTH-1) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL TMP_RAM: RAM_TYPE := (

         0 => x"3C080000", -- lui $t0, 0000
         1 => x"2508082C", -- addiu $t0, $t0, 2092
         2 => x"3C090000", -- lui $t1, 0000
         3 => x"25290840", -- addiu $t1, $t1, 2112
         4 => x"11090003", -- beq $t0, $t1, 3
         5 => x"25080004", -- addiu $t0, $t0, 4
         6 => x"08000004", -- j 4
         7 => x"AD00FFFC", -- sw $zero, -4(t0)
         8 => x"00000821", -- addu $at, $zero, $zero
         9 => x"00001021", -- addu $v0, $zero, $zero
        10 => x"00001821", -- addu $v1, $zero, $zero
        11 => x"00002021", -- addu $a0, $zero, $zero
        12 => x"00002821", -- addu $a1, $zero, $zero
        13 => x"00003021", -- addu $a2, $zero, $zero
        14 => x"00003821", -- addu $a3, $zero, $zero
        15 => x"00004021", -- addu $t0, $zero, $zero
        16 => x"00004821", -- addu $t1, $zero, $zero
        17 => x"00005021", -- addu $t2, $zero, $zero
        18 => x"00005821", -- addu $t3, $zero, $zero
        19 => x"00006021", -- addu $t4, $zero, $zero
        20 => x"00006821", -- addu $t5, $zero, $zero
        21 => x"00007021", -- addu $t6, $zero, $zero
        22 => x"00007821", -- addu $t7, $zero, $zero
        23 => x"00008021", -- addu $s0, $zero, $zero
        24 => x"00008821", -- addu $s1, $zero, $zero
        25 => x"00009021", -- addu $s2, $zero, $zero
        26 => x"00009821", -- addu $s3, $zero, $zero
        27 => x"0000A021", -- addu $s4, $zero, $zero
        28 => x"0000A821", -- addu $s5, $zero, $zero
        29 => x"0000B021", -- addu $s6, $zero, $zero
        30 => x"0000B821", -- addu $s7, $zero, $zero
        31 => x"0000C021", -- addu $t8, $zero, $zero
        32 => x"0000C821", -- addu $t9, $zero, $zero
        33 => x"0000D021", -- addu $k0, $zero, $zero
        34 => x"0000D821", -- addu $k1, $zero, $zero
        35 => x"0000E021", -- addu $gp, $zero, $zero
        36 => x"0000F821", -- addu $ra, $zero, $zero
        37 => x"3C1D0000", -- lui $sp, 0000
        38 => x"27BD0FF8", -- addiu $sp, $sp, 4088
        39 => x"0C0001D9", -- jal 473
        40 => x"03A0F021", -- addu $fp, $sp, $zero
        41 => x"08000029", -- j 41
        42 => x"00000000", -- nop
        43 => x"27BDFE90", -- addiu $sp, $sp, -368
        44 => x"AFBE016C", -- sw $fp, 364(sp)
        45 => x"03A0F021", -- addu $fp, $sp, $zero
        46 => x"AFC40170", -- sw $a0, 368(fp)
        47 => x"AFC00000", -- sw $zero, 0(fp)
        48 => x"08000067", -- j 103
        49 => x"00000000", -- nop
        50 => x"8FC50000", -- lw $a1, 0(fp)
        51 => x"8FC20000", -- lw $v0, 0(fp)
        52 => x"00000000", -- nop
        53 => x"00021080", -- sll $v0, $v0, 4
        54 => x"00401821", -- addu $v1, $v0, $zero
        55 => x"8FC20170", -- lw $v0, 368(fp)
        56 => x"00000000", -- nop
        57 => x"00431021", -- addu $v0, $v0, $v1
        58 => x"90420000", -- lbu $v0, 0(v0)
        59 => x"00000000", -- nop
        60 => x"00022600", -- sll $a0, $v0, 16
        61 => x"8FC20000", -- lw $v0, 0(fp)
        62 => x"00000000", -- nop
        63 => x"00021080", -- sll $v0, $v0, 4
        64 => x"24430001", -- addiu $v1, $v0, 1
        65 => x"8FC20170", -- lw $v0, 368(fp)
        66 => x"00000000", -- nop
        67 => x"00431021", -- addu $v0, $v0, $v1
        68 => x"90420000", -- lbu $v0, 0(v0)
        69 => x"00000000", -- nop
        70 => x"00021400", -- sll $v0, $v0, 0
        71 => x"00822025", -- or $a0, $a0, $v0
        72 => x"8FC20000", -- lw $v0, 0(fp)
        73 => x"00000000", -- nop
        74 => x"00021040", -- sll $v0, $v0, 2
        75 => x"24420001", -- addiu $v0, $v0, 1
        76 => x"00021040", -- sll $v0, $v0, 2
        77 => x"00401821", -- addu $v1, $v0, $zero
        78 => x"8FC20170", -- lw $v0, 368(fp)
        79 => x"00000000", -- nop
        80 => x"00431021", -- addu $v0, $v0, $v1
        81 => x"90420000", -- lbu $v0, 0(v0)
        82 => x"00000000", -- nop
        83 => x"00021200", -- sll $v0, $v0, 16
        84 => x"00822025", -- or $a0, $a0, $v0
        85 => x"8FC20000", -- lw $v0, 0(fp)
        86 => x"00000000", -- nop
        87 => x"00021080", -- sll $v0, $v0, 4
        88 => x"24430003", -- addiu $v1, $v0, 3
        89 => x"8FC20170", -- lw $v0, 368(fp)
        90 => x"00000000", -- nop
        91 => x"00431021", -- addu $v0, $v0, $v1
        92 => x"90420000", -- lbu $v0, 0(v0)
        93 => x"00000000", -- nop
        94 => x"00821025", -- or $v0, $a0, $v0
        95 => x"00401821", -- addu $v1, $v0, $zero
        96 => x"00051080", -- sll $v0, $a1, 4
        97 => x"03C21021", -- addu $v0, $fp, $v0
        98 => x"AC430024", -- sw $v1, 36(v0)
        99 => x"8FC20000", -- lw $v0, 0(fp)
       100 => x"00000000", -- nop
       101 => x"24420001", -- addiu $v0, $v0, 1
       102 => x"AFC20000", -- sw $v0, 0(fp)
       103 => x"8FC20000", -- lw $v0, 0(fp)
       104 => x"00000000", -- nop
       105 => x"28420010", -- slti $v0, $v0, 16
       106 => x"1440FFC7", -- bne $v0, $zero, -57
       107 => x"00000000", -- nop
       108 => x"08000097", -- j 151
       109 => x"00000000", -- nop
       110 => x"8FC50000", -- lw $a1, 0(fp)
       111 => x"8FC20000", -- lw $v0, 0(fp)
       112 => x"00000000", -- nop
       113 => x"2442FFFD", -- addiu $v0, $v0, -3
       114 => x"00021080", -- sll $v0, $v0, 4
       115 => x"03C21021", -- addu $v0, $fp, $v0
       116 => x"8C430024", -- lw $v1, 36(v0)
       117 => x"8FC20000", -- lw $v0, 0(fp)
       118 => x"00000000", -- nop
       119 => x"2442FFF8", -- addiu $v0, $v0, -8
       120 => x"00021080", -- sll $v0, $v0, 4
       121 => x"03C21021", -- addu $v0, $fp, $v0
       122 => x"8C420024", -- lw $v0, 36(v0)
       123 => x"00000000", -- nop
       124 => x"00621826", -- xor $v1, $v1, $v0
       125 => x"8FC20000", -- lw $v0, 0(fp)
       126 => x"00000000", -- nop
       127 => x"2442FFF2", -- addiu $v0, $v0, -14
       128 => x"00021080", -- sll $v0, $v0, 4
       129 => x"03C21021", -- addu $v0, $fp, $v0
       130 => x"8C420024", -- lw $v0, 36(v0)
       131 => x"00000000", -- nop
       132 => x"00621826", -- xor $v1, $v1, $v0
       133 => x"8FC20000", -- lw $v0, 0(fp)
       134 => x"00000000", -- nop
       135 => x"2442FFF0", -- addiu $v0, $v0, -16
       136 => x"00021080", -- sll $v0, $v0, 4
       137 => x"03C21021", -- addu $v0, $fp, $v0
       138 => x"8C420024", -- lw $v0, 36(v0)
       139 => x"00000000", -- nop
       140 => x"00621026", -- xor $v0, $v1, $v0
       141 => x"000227C2", -- srl $a0, $v0, 30
       142 => x"00021840", -- sll $v1, $v0, 2
       143 => x"00641825", -- or $v1, $v1, $a0
       144 => x"00051080", -- sll $v0, $a1, 4
       145 => x"03C21021", -- addu $v0, $fp, $v0
       146 => x"AC430024", -- sw $v1, 36(v0)
       147 => x"8FC20000", -- lw $v0, 0(fp)
       148 => x"00000000", -- nop
       149 => x"24420001", -- addiu $v0, $v0, 1
       150 => x"AFC20000", -- sw $v0, 0(fp)
       151 => x"8FC20000", -- lw $v0, 0(fp)
       152 => x"00000000", -- nop
       153 => x"28420050", -- slti $v0, $v0, 80
       154 => x"1440FFD3", -- bne $v0, $zero, -45
       155 => x"00000000", -- nop
       156 => x"8F820834", -- lw $v0, 2100(gp)
       157 => x"00000000", -- nop
       158 => x"AFC20020", -- sw $v0, 32(fp)
       159 => x"8F82082C", -- lw $v0, 2092(gp)
       160 => x"00000000", -- nop
       161 => x"AFC2001C", -- sw $v0, 28(fp)
       162 => x"8F820830", -- lw $v0, 2096(gp)
       163 => x"00000000", -- nop
       164 => x"AFC20018", -- sw $v0, 24(fp)
       165 => x"8F82083C", -- lw $v0, 2108(gp)
       166 => x"00000000", -- nop
       167 => x"AFC20014", -- sw $v0, 20(fp)
       168 => x"8F820838", -- lw $v0, 2104(gp)
       169 => x"00000000", -- nop
       170 => x"AFC20010", -- sw $v0, 16(fp)
       171 => x"AFC00000", -- sw $zero, 0(fp)
       172 => x"08000124", -- j 292
       173 => x"00000000", -- nop
       174 => x"8FC20000", -- lw $v0, 0(fp)
       175 => x"00000000", -- nop
       176 => x"28420014", -- slti $v0, $v0, 20
       177 => x"10400012", -- beq $v0, $zero, 18
       178 => x"00000000", -- nop
       179 => x"8FC3001C", -- lw $v1, 28(fp)
       180 => x"8FC20018", -- lw $v0, 24(fp)
       181 => x"00000000", -- nop
       182 => x"00622024", -- and $a0, $v1, $v0
       183 => x"8FC2001C", -- lw $v0, 28(fp)
       184 => x"00000000", -- nop
       185 => x"00021827", -- nor $v1, $zero, $v0
       186 => x"8FC20014", -- lw $v0, 20(fp)
       187 => x"00000000", -- nop
       188 => x"00621024", -- and $v0, $v1, $v0
       189 => x"00821025", -- or $v0, $a0, $v0
       190 => x"AFC2000C", -- sw $v0, 12(fp)
       191 => x"3C025A82", -- lui $v0, 5a82
       192 => x"34427999", -- ori $v0, $v0, 7999
       193 => x"AFC20008", -- sw $v0, 8(fp)
       194 => x"080000F8", -- j 248
       195 => x"00000000", -- nop
       196 => x"8FC20000", -- lw $v0, 0(fp)
       197 => x"00000000", -- nop
       198 => x"28420028", -- slti $v0, $v0, 40
       199 => x"1040000E", -- beq $v0, $zero, 14
       200 => x"00000000", -- nop
       201 => x"8FC3001C", -- lw $v1, 28(fp)
       202 => x"8FC20018", -- lw $v0, 24(fp)
       203 => x"00000000", -- nop
       204 => x"00621826", -- xor $v1, $v1, $v0
       205 => x"8FC20014", -- lw $v0, 20(fp)
       206 => x"00000000", -- nop
       207 => x"00621026", -- xor $v0, $v1, $v0
       208 => x"AFC2000C", -- sw $v0, 12(fp)
       209 => x"3C026ED9", -- lui $v0, 6ed9
       210 => x"3442EBA1", -- ori $v0, $v0, eba1
       211 => x"AFC20008", -- sw $v0, 8(fp)
       212 => x"080000F8", -- j 248
       213 => x"00000000", -- nop
       214 => x"8FC20000", -- lw $v0, 0(fp)
       215 => x"00000000", -- nop
       216 => x"2842003C", -- slti $v0, $v0, 60
       217 => x"10400013", -- beq $v0, $zero, 19
       218 => x"00000000", -- nop
       219 => x"8FC30018", -- lw $v1, 24(fp)
       220 => x"8FC20014", -- lw $v0, 20(fp)
       221 => x"00000000", -- nop
       222 => x"00621825", -- or $v1, $v1, $v0
       223 => x"8FC2001C", -- lw $v0, 28(fp)
       224 => x"00000000", -- nop
       225 => x"00622024", -- and $a0, $v1, $v0
       226 => x"8FC30018", -- lw $v1, 24(fp)
       227 => x"8FC20014", -- lw $v0, 20(fp)
       228 => x"00000000", -- nop
       229 => x"00621024", -- and $v0, $v1, $v0
       230 => x"00821025", -- or $v0, $a0, $v0
       231 => x"AFC2000C", -- sw $v0, 12(fp)
       232 => x"3C028F1B", -- lui $v0, 8f1b
       233 => x"3442BCDC", -- ori $v0, $v0, bcdc
       234 => x"AFC20008", -- sw $v0, 8(fp)
       235 => x"080000F8", -- j 248
       236 => x"00000000", -- nop
       237 => x"8FC3001C", -- lw $v1, 28(fp)
       238 => x"8FC20018", -- lw $v0, 24(fp)
       239 => x"00000000", -- nop
       240 => x"00621826", -- xor $v1, $v1, $v0
       241 => x"8FC20014", -- lw $v0, 20(fp)
       242 => x"00000000", -- nop
       243 => x"00621026", -- xor $v0, $v1, $v0
       244 => x"AFC2000C", -- sw $v0, 12(fp)
       245 => x"3C02CA62", -- lui $v0, ca62
       246 => x"3442C1D6", -- ori $v0, $v0, c1d6
       247 => x"AFC20008", -- sw $v0, 8(fp)
       248 => x"8FC20020", -- lw $v0, 32(fp)
       249 => x"00000000", -- nop
       250 => x"00021EC2", -- srl $v1, $v0, 22
       251 => x"00021140", -- sll $v0, $v0, 10
       252 => x"00431025", -- or $v0, $v0, $v1
       253 => x"8FC3000C", -- lw $v1, 12(fp)
       254 => x"00000000", -- nop
       255 => x"00431821", -- addu $v1, $v0, $v1
       256 => x"8FC20010", -- lw $v0, 16(fp)
       257 => x"00000000", -- nop
       258 => x"00621821", -- addu $v1, $v1, $v0
       259 => x"8FC20008", -- lw $v0, 8(fp)
       260 => x"00000000", -- nop
       261 => x"00621821", -- addu $v1, $v1, $v0
       262 => x"8FC20000", -- lw $v0, 0(fp)
       263 => x"00000000", -- nop
       264 => x"00021080", -- sll $v0, $v0, 4
       265 => x"03C21021", -- addu $v0, $fp, $v0
       266 => x"8C420024", -- lw $v0, 36(v0)
       267 => x"00000000", -- nop
       268 => x"00621021", -- addu $v0, $v1, $v0
       269 => x"AFC20004", -- sw $v0, 4(fp)
       270 => x"8FC20014", -- lw $v0, 20(fp)
       271 => x"00000000", -- nop
       272 => x"AFC20010", -- sw $v0, 16(fp)
       273 => x"8FC20018", -- lw $v0, 24(fp)
       274 => x"00000000", -- nop
       275 => x"AFC20014", -- sw $v0, 20(fp)
       276 => x"8FC2001C", -- lw $v0, 28(fp)
       277 => x"00000000", -- nop
       278 => x"00021882", -- srl $v1, $v0, 4
       279 => x"00021780", -- sll $v0, $v0, 28
       280 => x"00621025", -- or $v0, $v1, $v0
       281 => x"AFC20018", -- sw $v0, 24(fp)
       282 => x"8FC20020", -- lw $v0, 32(fp)
       283 => x"00000000", -- nop
       284 => x"AFC2001C", -- sw $v0, 28(fp)
       285 => x"8FC20004", -- lw $v0, 4(fp)
       286 => x"00000000", -- nop
       287 => x"AFC20020", -- sw $v0, 32(fp)
       288 => x"8FC20000", -- lw $v0, 0(fp)
       289 => x"00000000", -- nop
       290 => x"24420001", -- addiu $v0, $v0, 1
       291 => x"AFC20000", -- sw $v0, 0(fp)
       292 => x"8FC20000", -- lw $v0, 0(fp)
       293 => x"00000000", -- nop
       294 => x"28420050", -- slti $v0, $v0, 80
       295 => x"1440FF86", -- bne $v0, $zero, -122
       296 => x"00000000", -- nop
       297 => x"8F830834", -- lw $v1, 2100(gp)
       298 => x"8FC20020", -- lw $v0, 32(fp)
       299 => x"00000000", -- nop
       300 => x"00621021", -- addu $v0, $v1, $v0
       301 => x"AF820834", -- sw $v0, 2100(gp)
       302 => x"8F83082C", -- lw $v1, 2092(gp)
       303 => x"8FC2001C", -- lw $v0, 28(fp)
       304 => x"00000000", -- nop
       305 => x"00621021", -- addu $v0, $v1, $v0
       306 => x"AF82082C", -- sw $v0, 2092(gp)
       307 => x"8F830830", -- lw $v1, 2096(gp)
       308 => x"8FC20018", -- lw $v0, 24(fp)
       309 => x"00000000", -- nop
       310 => x"00621021", -- addu $v0, $v1, $v0
       311 => x"AF820830", -- sw $v0, 2096(gp)
       312 => x"8F83083C", -- lw $v1, 2108(gp)
       313 => x"8FC20014", -- lw $v0, 20(fp)
       314 => x"00000000", -- nop
       315 => x"00621021", -- addu $v0, $v1, $v0
       316 => x"AF82083C", -- sw $v0, 2108(gp)
       317 => x"8F830838", -- lw $v1, 2104(gp)
       318 => x"8FC20010", -- lw $v0, 16(fp)
       319 => x"00000000", -- nop
       320 => x"00621021", -- addu $v0, $v1, $v0
       321 => x"AF820838", -- sw $v0, 2104(gp)
       322 => x"03C0E821", -- addu $sp, $fp, $zero
       323 => x"8FBE016C", -- lw $fp, 364(sp)
       324 => x"27BD0170", -- addiu $sp, $sp, 368
       325 => x"03E00008", -- jr $ra
       326 => x"00000000", -- nop
       327 => x"27BDFF98", -- addiu $sp, $sp, -104
       328 => x"AFBF0064", -- sw $ra, 100(sp)
       329 => x"AFBE0060", -- sw $fp, 96(sp)
       330 => x"03A0F021", -- addu $fp, $sp, $zero
       331 => x"AFC40068", -- sw $a0, 104(fp)
       332 => x"AFC5006C", -- sw $a1, 108(fp)
       333 => x"3C026745", -- lui $v0, 6745
       334 => x"34422301", -- ori $v0, $v0, 2301
       335 => x"AF820834", -- sw $v0, 2100(gp)
       336 => x"3C02EFCD", -- lui $v0, efcd
       337 => x"3442AB89", -- ori $v0, $v0, ab89
       338 => x"AF82082C", -- sw $v0, 2092(gp)
       339 => x"3C0298BA", -- lui $v0, 98ba
       340 => x"3442DCFE", -- ori $v0, $v0, dcfe
       341 => x"AF820830", -- sw $v0, 2096(gp)
       342 => x"3C021032", -- lui $v0, 1032
       343 => x"34425476", -- ori $v0, $v0, 5476
       344 => x"AF82083C", -- sw $v0, 2108(gp)
       345 => x"3C02C3D2", -- lui $v0, c3d2
       346 => x"3442E1F0", -- ori $v0, $v0, e1f0
       347 => x"AF820838", -- sw $v0, 2104(gp)
       348 => x"8FC2006C", -- lw $v0, 108(fp)
       349 => x"00000000", -- nop
       350 => x"AFC20010", -- sw $v0, 16(fp)
       351 => x"0800016C", -- j 364
       352 => x"00000000", -- nop
       353 => x"8FC40068", -- lw $a0, 104(fp)
       354 => x"0C00002B", -- jal 43
       355 => x"00000000", -- nop
       356 => x"8FC20068", -- lw $v0, 104(fp)
       357 => x"00000000", -- nop
       358 => x"24420040", -- addiu $v0, $v0, 64
       359 => x"AFC20068", -- sw $v0, 104(fp)
       360 => x"8FC20010", -- lw $v0, 16(fp)
       361 => x"00000000", -- nop
       362 => x"2442FFC0", -- addiu $v0, $v0, -64
       363 => x"AFC20010", -- sw $v0, 16(fp)
       364 => x"8FC20010", -- lw $v0, 16(fp)
       365 => x"00000000", -- nop
       366 => x"28420040", -- slti $v0, $v0, 64
       367 => x"1040FFF1", -- beq $v0, $zero, -15
       368 => x"00000000", -- nop
       369 => x"AFC00014", -- sw $zero, 20(fp)
       370 => x"08000192", -- j 402
       371 => x"00000000", -- nop
       372 => x"8FC20014", -- lw $v0, 20(fp)
       373 => x"00000000", -- nop
       374 => x"AFC2005C", -- sw $v0, 92(fp)
       375 => x"8FC20014", -- lw $v0, 20(fp)
       376 => x"8FC30010", -- lw $v1, 16(fp)
       377 => x"00000000", -- nop
       378 => x"0043102A", -- slt $v0, $v0, $v1
       379 => x"1040000A", -- beq $v0, $zero, 10
       380 => x"00000000", -- nop
       381 => x"8FC20014", -- lw $v0, 20(fp)
       382 => x"8FC30068", -- lw $v1, 104(fp)
       383 => x"00000000", -- nop
       384 => x"00621021", -- addu $v0, $v1, $v0
       385 => x"90420000", -- lbu $v0, 0(v0)
       386 => x"00000000", -- nop
       387 => x"AFC20058", -- sw $v0, 88(fp)
       388 => x"08000187", -- j 391
       389 => x"00000000", -- nop
       390 => x"AFC00058", -- sw $zero, 88(fp)
       391 => x"27C20010", -- addiu $v0, $fp, 16
       392 => x"8FC3005C", -- lw $v1, 92(fp)
       393 => x"00000000", -- nop
       394 => x"00431021", -- addu $v0, $v0, $v1
       395 => x"8FC30058", -- lw $v1, 88(fp)
       396 => x"00000000", -- nop
       397 => x"A0430008", -- sb $v1, 8(v0)
       398 => x"8FC20014", -- lw $v0, 20(fp)
       399 => x"00000000", -- nop
       400 => x"24420001", -- addiu $v0, $v0, 1
       401 => x"AFC20014", -- sw $v0, 20(fp)
       402 => x"8FC20014", -- lw $v0, 20(fp)
       403 => x"00000000", -- nop
       404 => x"28420040", -- slti $v0, $v0, 64
       405 => x"1440FFDE", -- bne $v0, $zero, -34
       406 => x"00000000", -- nop
       407 => x"8FC30010", -- lw $v1, 16(fp)
       408 => x"27C20010", -- addiu $v0, $fp, 16
       409 => x"00431821", -- addu $v1, $v0, $v1
       410 => x"2402FF80", -- addiu $v0, $zero, -128
       411 => x"A0620008", -- sb $v0, 8(v1)
       412 => x"8FC20010", -- lw $v0, 16(fp)
       413 => x"00000000", -- nop
       414 => x"28420038", -- slti $v0, $v0, 56
       415 => x"14400015", -- bne $v0, $zero, 21
       416 => x"00000000", -- nop
       417 => x"27C20018", -- addiu $v0, $fp, 24
       418 => x"00402021", -- addu $a0, $v0, $zero
       419 => x"0C00002B", -- jal 43
       420 => x"00000000", -- nop
       421 => x"AFC00014", -- sw $zero, 20(fp)
       422 => x"080001B0", -- j 432
       423 => x"00000000", -- nop
       424 => x"8FC30014", -- lw $v1, 20(fp)
       425 => x"27C20010", -- addiu $v0, $fp, 16
       426 => x"00431021", -- addu $v0, $v0, $v1
       427 => x"A0400008", -- sb $zero, 8(v0)
       428 => x"8FC20014", -- lw $v0, 20(fp)
       429 => x"00000000", -- nop
       430 => x"24420001", -- addiu $v0, $v0, 1
       431 => x"AFC20014", -- sw $v0, 20(fp)
       432 => x"8FC20014", -- lw $v0, 20(fp)
       433 => x"00000000", -- nop
       434 => x"2842003B", -- slti $v0, $v0, 59
       435 => x"1440FFF4", -- bne $v0, $zero, -12
       436 => x"00000000", -- nop
       437 => x"8FC2006C", -- lw $v0, 108(fp)
       438 => x"00000000", -- nop
       439 => x"00021742", -- srl $v0, $v0, 26
       440 => x"304200FF", -- andi $v0, $v0, 00ff
       441 => x"A3C20053", -- sb $v0, 83(fp)
       442 => x"8FC2006C", -- lw $v0, 108(fp)
       443 => x"00000000", -- nop
       444 => x"00021542", -- srl $v0, $v0, 10
       445 => x"304200FF", -- andi $v0, $v0, 00ff
       446 => x"A3C20054", -- sb $v0, 84(fp)
       447 => x"8FC2006C", -- lw $v0, 108(fp)
       448 => x"00000000", -- nop
       449 => x"00021342", -- srl $v0, $v0, 26
       450 => x"304200FF", -- andi $v0, $v0, 00ff
       451 => x"A3C20055", -- sb $v0, 85(fp)
       452 => x"8FC2006C", -- lw $v0, 108(fp)
       453 => x"00000000", -- nop
       454 => x"00021142", -- srl $v0, $v0, 10
       455 => x"304200FF", -- andi $v0, $v0, 00ff
       456 => x"A3C20056", -- sb $v0, 86(fp)
       457 => x"8FC2006C", -- lw $v0, 108(fp)
       458 => x"00000000", -- nop
       459 => x"304200FF", -- andi $v0, $v0, 00ff
       460 => x"000210C0", -- sll $v0, $v0, 6
       461 => x"304200FF", -- andi $v0, $v0, 00ff
       462 => x"A3C20057", -- sb $v0, 87(fp)
       463 => x"27C20018", -- addiu $v0, $fp, 24
       464 => x"00402021", -- addu $a0, $v0, $zero
       465 => x"0C00002B", -- jal 43
       466 => x"00000000", -- nop
       467 => x"03C0E821", -- addu $sp, $fp, $zero
       468 => x"8FBF0064", -- lw $ra, 100(sp)
       469 => x"8FBE0060", -- lw $fp, 96(sp)
       470 => x"27BD0068", -- addiu $sp, $sp, 104
       471 => x"03E00008", -- jr $ra
       472 => x"00000000", -- nop
       473 => x"27BDFFE8", -- addiu $sp, $sp, -24
       474 => x"AFBF0014", -- sw $ra, 20(sp)
       475 => x"AFBE0010", -- sw $fp, 16(sp)
       476 => x"03A0F021", -- addu $fp, $sp, $zero
       477 => x"3C020000", -- lui $v0, 0000
       478 => x"24420800", -- addiu $v0, $v0, 2048
       479 => x"00402021", -- addu $a0, $v0, $zero
       480 => x"2405002B", -- addiu $a1, $zero, 43
       481 => x"0C000147", -- jal 327
       482 => x"00000000", -- nop
       483 => x"00001021", -- addu $v0, $zero, $zero
       484 => x"03C0E821", -- addu $sp, $fp, $zero
       485 => x"8FBF0014", -- lw $ra, 20(sp)
       486 => x"8FBE0010", -- lw $fp, 16(sp)
       487 => x"27BD0018", -- addiu $sp, $sp, 24
       488 => x"03E00008", -- jr $ra
       489 => x"00000000", -- nop
       490 => x"00000000", -- nop
       491 => x"00000000", -- nop
       492 => x"00000000", -- nop
       493 => x"00000000", -- nop
       494 => x"00000000", -- nop
       495 => x"00000000", -- nop
       496 => x"00000000", -- nop
       497 => x"00000000", -- nop
       498 => x"00000000", -- nop
       499 => x"00000000", -- nop
       500 => x"00000000", -- nop
       501 => x"00000000", -- nop
       502 => x"00000000", -- nop
       503 => x"00000000", -- nop
       504 => x"00000000", -- nop
       505 => x"00000000", -- nop
       506 => x"00000000", -- nop
       507 => x"00000000", -- nop
       508 => x"00000000", -- nop
       509 => x"00000000", -- nop
       510 => x"00000000", -- nop
       511 => x"00000000"  -- nop
    );

BEGIN

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF R='1' THEN
                DATA_OUT <= TMP_RAM(CONV_INTEGER(UNSIGNED(RADDR(ADDR-1 DOWNTO 2))));
            ELSE
                DATA_OUT <= (DATA_OUT'RANGE => 'Z');
            END IF;
        END IF;
    END IF;
    END PROCESS;

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF W='1' THEN
                TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2)))) <= DATA_IN;
            END IF;
        END IF;
    END IF;
    END PROCESS;

END BEHAV_CODE;

ARCHITECTURE BEHAV_DATA OF SRAM IS

    TYPE RAM_TYPE IS ARRAY (0 TO DEPTH-1) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL IBYTE0:     STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL IBYTE1:     STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL IBYTE2:     STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL IBYTE3:     STD_LOGIC_VECTOR(7 DOWNTO 0);

    SIGNAL OBYTE:      STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL OHALF:      STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SBYTE:      STD_LOGIC_VECTOR(23 DOWNTO 0);
    SIGNAL SHALF:      STD_LOGIC_VECTOR(15 DOWNTO 0);

    SIGNAL RWORD:      STD_LOGIC_VECTOR(31 DOWNTO 0):= x"00000000";

    SIGNAL RADDR2:     STD_LOGIC_VECTOR(1 DOWNTO 0):= "00";
    SIGNAL MODE2:      STD_LOGIC_VECTOR(2 DOWNTO 0):= "000";
    SIGNAL ISSIGNED2:  STD_LOGIC:= '0';

    SIGNAL W0:         STD_LOGIC;
    SIGNAL W1:         STD_LOGIC;
    SIGNAL W2:         STD_LOGIC;
    SIGNAL W3:         STD_LOGIC;

    SIGNAL TMP_RAM: RAM_TYPE := (

         0 => x"54686520",
         1 => x"71756963",
         2 => x"6B206272",
         3 => x"6F776E20",
         4 => x"666F7820",
         5 => x"6A756D70",
         6 => x"73206F76",
         7 => x"65722074",
         8 => x"6865206C",
         9 => x"617A7920",
        10 => x"646F6700",
        11 => x"55555555",
        12 => x"55555555",
        13 => x"55555555",
        14 => x"55555555",
        15 => x"55555555",
        16 => x"55555555",
        17 => x"55555555",
        18 => x"55555555",
        19 => x"55555555",
        20 => x"55555555",
        21 => x"55555555",
        22 => x"55555555",
        23 => x"55555555",
        24 => x"55555555",
        25 => x"55555555",
        26 => x"55555555",
        27 => x"55555555",
        28 => x"55555555",
        29 => x"55555555",
        30 => x"55555555",
        31 => x"55555555",
        32 => x"55555555",
        33 => x"55555555",
        34 => x"55555555",
        35 => x"55555555",
        36 => x"55555555",
        37 => x"55555555",
        38 => x"55555555",
        39 => x"55555555",
        40 => x"55555555",
        41 => x"55555555",
        42 => x"55555555",
        43 => x"55555555",
        44 => x"55555555",
        45 => x"55555555",
        46 => x"55555555",
        47 => x"55555555",
        48 => x"55555555",
        49 => x"55555555",
        50 => x"55555555",
        51 => x"55555555",
        52 => x"55555555",
        53 => x"55555555",
        54 => x"55555555",
        55 => x"55555555",
        56 => x"55555555",
        57 => x"55555555",
        58 => x"55555555",
        59 => x"55555555",
        60 => x"55555555",
        61 => x"55555555",
        62 => x"55555555",
        63 => x"55555555",
        64 => x"55555555",
        65 => x"55555555",
        66 => x"55555555",
        67 => x"55555555",
        68 => x"55555555",
        69 => x"55555555",
        70 => x"55555555",
        71 => x"55555555",
        72 => x"55555555",
        73 => x"55555555",
        74 => x"55555555",
        75 => x"55555555",
        76 => x"55555555",
        77 => x"55555555",
        78 => x"55555555",
        79 => x"55555555",
        80 => x"55555555",
        81 => x"55555555",
        82 => x"55555555",
        83 => x"55555555",
        84 => x"55555555",
        85 => x"55555555",
        86 => x"55555555",
        87 => x"55555555",
        88 => x"55555555",
        89 => x"55555555",
        90 => x"55555555",
        91 => x"55555555",
        92 => x"55555555",
        93 => x"55555555",
        94 => x"55555555",
        95 => x"55555555",
        96 => x"55555555",
        97 => x"55555555",
        98 => x"55555555",
        99 => x"55555555",
       100 => x"55555555",
       101 => x"55555555",
       102 => x"55555555",
       103 => x"55555555",
       104 => x"55555555",
       105 => x"55555555",
       106 => x"55555555",
       107 => x"55555555",
       108 => x"55555555",
       109 => x"55555555",
       110 => x"55555555",
       111 => x"55555555",
       112 => x"55555555",
       113 => x"55555555",
       114 => x"55555555",
       115 => x"55555555",
       116 => x"55555555",
       117 => x"55555555",
       118 => x"55555555",
       119 => x"55555555",
       120 => x"55555555",
       121 => x"55555555",
       122 => x"55555555",
       123 => x"55555555",
       124 => x"55555555",
       125 => x"55555555",
       126 => x"55555555",
       127 => x"55555555",
       128 => x"55555555",
       129 => x"55555555",
       130 => x"55555555",
       131 => x"55555555",
       132 => x"55555555",
       133 => x"55555555",
       134 => x"55555555",
       135 => x"55555555",
       136 => x"55555555",
       137 => x"55555555",
       138 => x"55555555",
       139 => x"55555555",
       140 => x"55555555",
       141 => x"55555555",
       142 => x"55555555",
       143 => x"55555555",
       144 => x"55555555",
       145 => x"55555555",
       146 => x"55555555",
       147 => x"55555555",
       148 => x"55555555",
       149 => x"55555555",
       150 => x"55555555",
       151 => x"55555555",
       152 => x"55555555",
       153 => x"55555555",
       154 => x"55555555",
       155 => x"55555555",
       156 => x"55555555",
       157 => x"55555555",
       158 => x"55555555",
       159 => x"55555555",
       160 => x"55555555",
       161 => x"55555555",
       162 => x"55555555",
       163 => x"55555555",
       164 => x"55555555",
       165 => x"55555555",
       166 => x"55555555",
       167 => x"55555555",
       168 => x"55555555",
       169 => x"55555555",
       170 => x"55555555",
       171 => x"55555555",
       172 => x"55555555",
       173 => x"55555555",
       174 => x"55555555",
       175 => x"55555555",
       176 => x"55555555",
       177 => x"55555555",
       178 => x"55555555",
       179 => x"55555555",
       180 => x"55555555",
       181 => x"55555555",
       182 => x"55555555",
       183 => x"55555555",
       184 => x"55555555",
       185 => x"55555555",
       186 => x"55555555",
       187 => x"55555555",
       188 => x"55555555",
       189 => x"55555555",
       190 => x"55555555",
       191 => x"55555555",
       192 => x"55555555",
       193 => x"55555555",
       194 => x"55555555",
       195 => x"55555555",
       196 => x"55555555",
       197 => x"55555555",
       198 => x"55555555",
       199 => x"55555555",
       200 => x"55555555",
       201 => x"55555555",
       202 => x"55555555",
       203 => x"55555555",
       204 => x"55555555",
       205 => x"55555555",
       206 => x"55555555",
       207 => x"55555555",
       208 => x"55555555",
       209 => x"55555555",
       210 => x"55555555",
       211 => x"55555555",
       212 => x"55555555",
       213 => x"55555555",
       214 => x"55555555",
       215 => x"55555555",
       216 => x"55555555",
       217 => x"55555555",
       218 => x"55555555",
       219 => x"55555555",
       220 => x"55555555",
       221 => x"55555555",
       222 => x"55555555",
       223 => x"55555555",
       224 => x"55555555",
       225 => x"55555555",
       226 => x"55555555",
       227 => x"55555555",
       228 => x"55555555",
       229 => x"55555555",
       230 => x"55555555",
       231 => x"55555555",
       232 => x"55555555",
       233 => x"55555555",
       234 => x"55555555",
       235 => x"55555555",
       236 => x"55555555",
       237 => x"55555555",
       238 => x"55555555",
       239 => x"55555555",
       240 => x"55555555",
       241 => x"55555555",
       242 => x"55555555",
       243 => x"55555555",
       244 => x"55555555",
       245 => x"55555555",
       246 => x"55555555",
       247 => x"55555555",
       248 => x"55555555",
       249 => x"55555555",
       250 => x"55555555",
       251 => x"55555555",
       252 => x"55555555",
       253 => x"55555555",
       254 => x"55555555",
       255 => x"55555555",
       256 => x"55555555",
       257 => x"55555555",
       258 => x"55555555",
       259 => x"55555555",
       260 => x"55555555",
       261 => x"55555555",
       262 => x"55555555",
       263 => x"55555555",
       264 => x"55555555",
       265 => x"55555555",
       266 => x"55555555",
       267 => x"55555555",
       268 => x"55555555",
       269 => x"55555555",
       270 => x"55555555",
       271 => x"55555555",
       272 => x"55555555",
       273 => x"55555555",
       274 => x"55555555",
       275 => x"55555555",
       276 => x"55555555",
       277 => x"55555555",
       278 => x"55555555",
       279 => x"55555555",
       280 => x"55555555",
       281 => x"55555555",
       282 => x"55555555",
       283 => x"55555555",
       284 => x"55555555",
       285 => x"55555555",
       286 => x"55555555",
       287 => x"55555555",
       288 => x"55555555",
       289 => x"55555555",
       290 => x"55555555",
       291 => x"55555555",
       292 => x"55555555",
       293 => x"55555555",
       294 => x"55555555",
       295 => x"55555555",
       296 => x"55555555",
       297 => x"55555555",
       298 => x"55555555",
       299 => x"55555555",
       300 => x"55555555",
       301 => x"55555555",
       302 => x"55555555",
       303 => x"55555555",
       304 => x"55555555",
       305 => x"55555555",
       306 => x"55555555",
       307 => x"55555555",
       308 => x"55555555",
       309 => x"55555555",
       310 => x"55555555",
       311 => x"55555555",
       312 => x"55555555",
       313 => x"55555555",
       314 => x"55555555",
       315 => x"55555555",
       316 => x"55555555",
       317 => x"55555555",
       318 => x"55555555",
       319 => x"55555555",
       320 => x"55555555",
       321 => x"55555555",
       322 => x"55555555",
       323 => x"55555555",
       324 => x"55555555",
       325 => x"55555555",
       326 => x"55555555",
       327 => x"55555555",
       328 => x"55555555",
       329 => x"55555555",
       330 => x"55555555",
       331 => x"55555555",
       332 => x"55555555",
       333 => x"55555555",
       334 => x"55555555",
       335 => x"55555555",
       336 => x"55555555",
       337 => x"55555555",
       338 => x"55555555",
       339 => x"55555555",
       340 => x"55555555",
       341 => x"55555555",
       342 => x"55555555",
       343 => x"55555555",
       344 => x"55555555",
       345 => x"55555555",
       346 => x"55555555",
       347 => x"55555555",
       348 => x"55555555",
       349 => x"55555555",
       350 => x"55555555",
       351 => x"55555555",
       352 => x"55555555",
       353 => x"55555555",
       354 => x"55555555",
       355 => x"55555555",
       356 => x"55555555",
       357 => x"55555555",
       358 => x"55555555",
       359 => x"55555555",
       360 => x"55555555",
       361 => x"55555555",
       362 => x"55555555",
       363 => x"55555555",
       364 => x"55555555",
       365 => x"55555555",
       366 => x"55555555",
       367 => x"55555555",
       368 => x"55555555",
       369 => x"55555555",
       370 => x"55555555",
       371 => x"55555555",
       372 => x"55555555",
       373 => x"55555555",
       374 => x"55555555",
       375 => x"55555555",
       376 => x"55555555",
       377 => x"55555555",
       378 => x"55555555",
       379 => x"55555555",
       380 => x"55555555",
       381 => x"55555555",
       382 => x"55555555",
       383 => x"55555555",
       384 => x"55555555",
       385 => x"55555555",
       386 => x"55555555",
       387 => x"55555555",
       388 => x"55555555",
       389 => x"55555555",
       390 => x"55555555",
       391 => x"55555555",
       392 => x"55555555",
       393 => x"55555555",
       394 => x"55555555",
       395 => x"55555555",
       396 => x"55555555",
       397 => x"55555555",
       398 => x"55555555",
       399 => x"55555555",
       400 => x"55555555",
       401 => x"55555555",
       402 => x"55555555",
       403 => x"55555555",
       404 => x"55555555",
       405 => x"55555555",
       406 => x"55555555",
       407 => x"55555555",
       408 => x"55555555",
       409 => x"55555555",
       410 => x"55555555",
       411 => x"55555555",
       412 => x"55555555",
       413 => x"55555555",
       414 => x"55555555",
       415 => x"55555555",
       416 => x"55555555",
       417 => x"55555555",
       418 => x"55555555",
       419 => x"55555555",
       420 => x"55555555",
       421 => x"55555555",
       422 => x"55555555",
       423 => x"55555555",
       424 => x"55555555",
       425 => x"55555555",
       426 => x"55555555",
       427 => x"55555555",
       428 => x"55555555",
       429 => x"55555555",
       430 => x"55555555",
       431 => x"55555555",
       432 => x"55555555",
       433 => x"55555555",
       434 => x"55555555",
       435 => x"55555555",
       436 => x"55555555",
       437 => x"55555555",
       438 => x"55555555",
       439 => x"55555555",
       440 => x"55555555",
       441 => x"55555555",
       442 => x"55555555",
       443 => x"55555555",
       444 => x"55555555",
       445 => x"55555555",
       446 => x"55555555",
       447 => x"55555555",
       448 => x"55555555",
       449 => x"55555555",
       450 => x"55555555",
       451 => x"55555555",
       452 => x"55555555",
       453 => x"55555555",
       454 => x"55555555",
       455 => x"55555555",
       456 => x"55555555",
       457 => x"55555555",
       458 => x"55555555",
       459 => x"55555555",
       460 => x"55555555",
       461 => x"55555555",
       462 => x"55555555",
       463 => x"55555555",
       464 => x"55555555",
       465 => x"55555555",
       466 => x"55555555",
       467 => x"55555555",
       468 => x"55555555",
       469 => x"55555555",
       470 => x"55555555",
       471 => x"55555555",
       472 => x"55555555",
       473 => x"55555555",
       474 => x"55555555",
       475 => x"55555555",
       476 => x"55555555",
       477 => x"55555555",
       478 => x"55555555",
       479 => x"55555555",
       480 => x"55555555",
       481 => x"55555555",
       482 => x"55555555",
       483 => x"55555555",
       484 => x"55555555",
       485 => x"55555555",
       486 => x"55555555",
       487 => x"55555555",
       488 => x"55555555",
       489 => x"55555555",
       490 => x"55555555",
       491 => x"55555555",
       492 => x"55555555",
       493 => x"55555555",
       494 => x"55555555",
       495 => x"55555555",
       496 => x"55555555",
       497 => x"55555555",
       498 => x"55555555",
       499 => x"55555555",
       500 => x"55555555",
       501 => x"55555555",
       502 => x"55555555",
       503 => x"55555555",
       504 => x"55555555",
       505 => x"55555555",
       506 => x"55555555",
       507 => x"55555555",
       508 => x"55555555",
       509 => x"55555555",
       510 => x"55555555",
       511 => x"55555555"
    );

BEGIN
    -- READ LOGIC
    OBYTE    <=      RWORD(31 DOWNTO 24) WHEN RADDR2(1 DOWNTO 0) = "00"
                ELSE RWORD(23 DOWNTO 16) WHEN RADDR2(1 DOWNTO 0) = "01"
                ELSE RWORD(15 DOWNTO  8) WHEN RADDR2(1 DOWNTO 0) = "10"
                ELSE RWORD( 7 DOWNTO  0);

    OHALF    <=      RWORD(31 DOWNTO 16) WHEN RADDR2(1 DOWNTO 0) = "00"
                ELSE RWORD(15 DOWNTO  0); -- THIS IS CASE "11", WE DON'T HANDLE THE OTHER CASES


    SBYTE    <=      x"FFFFFF" WHEN (OBYTE(7)  AND ISSIGNED2) = '1' ELSE x"000000";
    SHALF    <=      x"FFFF"   WHEN (OHALF(15) AND ISSIGNED2) = '1' ELSE x"0000";


    DATA_OUT <=      SBYTE & OBYTE WHEN MODE2(2) = '1'
                ELSE SHALF & OHALF WHEN MODE2(1) = '1'
                ELSE RWORD WHEN MODE2(0) = '1';

    -- WRITE LOGIC

    IBYTE0 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN(15 DOWNTO 8) WHEN MODE(1)='1' ELSE DATA_IN(31 DOWNTO  24);
    IBYTE1 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN( 7 DOWNTO 0) WHEN MODE(1)='1' ELSE DATA_IN(23 DOWNTO  16);
    IBYTE2 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN(15 DOWNTO 8) WHEN MODE(1)='1' ELSE DATA_IN(15 DOWNTO   8);
    IBYTE3 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN( 7 DOWNTO 0) WHEN MODE(1)='1' ELSE DATA_IN( 7 DOWNTO   0);

    W0 <= (   (MODE(2) AND NOT(WADDR(1) OR   WADDR(0)))  --B: "00"
           OR (MODE(1) AND NOT(WADDR(1)))                --H: "0x"
           OR  MODE(0)) AND W;                           --W: "Xx"
    W1 <= (   (MODE(2) AND NOT(WADDR(1)) AND WADDR(0))   --B: "01"
           OR (MODE(1) AND NOT(WADDR(1)))                --H: "0x"
           OR  MODE(0)) AND W;                           --W: "Xx"
    W2 <= (   (MODE(2) AND NOT(WADDR(0)) AND WADDR(1))   --B: "10"
           OR (MODE(1) AND     WADDR(1))                 --H: "1x"
           OR  MODE(0)) AND W;                           --W: "Xx"
    W3 <= (   (MODE(2) AND     WADDR(1) AND  WADDR(0))   --B: "11"
           OR (MODE(1) AND     WADDR(1))                 --H: "1x"
           OR  MODE(0)) AND W;                           --W: "Xx"

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        MODE2     <= MODE;
        ISSIGNED2 <= ISSIGNED;
        RADDR2 <= RADDR(1 DOWNTO 0);
    END IF;
    END PROCESS;

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF R='1' THEN
                RWORD <= TMP_RAM(CONV_INTEGER(UNSIGNED(RADDR(ADDR-1 DOWNTO 2))));
            ELSE
                RWORD <= (DATA_OUT'RANGE => 'Z');
            END IF;
        END IF;
    END IF;
    END PROCESS;

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF W='1' THEN
                IF W0 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(31 DOWNTO 24) <= IBYTE0;
                END IF;
                IF W1 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(23 DOWNTO 16) <= IBYTE1;
                END IF;
                IF W2 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(15 DOWNTO  8) <= IBYTE2;
                END IF;
                IF W3 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(7  DOWNTO  0) <= IBYTE3;
                END IF;
            END IF;
        END IF;
    END IF;
    END PROCESS;

END BEHAV_DATA;
