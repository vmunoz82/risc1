----------------------------------------------------------
--
-- 32 bits pipelined RISC processor
-- Copyright (c) 2010 Victor Munoz. All rights reserved.
-- derechos reservados, prohibida su reproduccion
--
-- Author: Victor Munoz
-- Contact: vmunoz@ingenieria-inversa.cl
--
----------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

----------------------------------------------------------

ENTITY SRAM IS
    GENERIC(
        ADDR:     INTEGER:= (9+2);
        DEPTH:    INTEGER:= 512
    );
    PORT(
        CLK:      IN  STD_LOGIC;
        ENABLE:   IN  STD_LOGIC;
        R:        IN  STD_LOGIC;
        W:        IN  STD_LOGIC;
        RADDR:    IN  STD_LOGIC_VECTOR(ADDR-1 DOWNTO 0);
        WADDR:    IN  STD_LOGIC_VECTOR(ADDR-1 DOWNTO 0);
        DATA_IN:  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
        MODE:     IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
        ISSIGNED: IN  STD_LOGIC;
        DATA_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0):= "00000000000000000000000000000000"
    );
END SRAM;

--------------------------------------------------------------

ARCHITECTURE BEHAV_CODE OF SRAM IS

    TYPE RAM_TYPE IS ARRAY (0 TO DEPTH-1) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL TMP_RAM: RAM_TYPE := (

         0 => x"3C080000", -- lui $t0, 0000
         1 => x"2508084C", -- addiu $t0, $t0, 2124
         2 => x"3C090000", -- lui $t1, 0000
         3 => x"25290854", -- addiu $t1, $t1, 2132
         4 => x"11090003", -- beq $t0, $t1, 3
         5 => x"25080004", -- addiu $t0, $t0, 4
         6 => x"08000004", -- j 4
         7 => x"AD00FFFC", -- sw $zero, -4(t0)
         8 => x"00000821", -- addu $at, $zero, $zero
         9 => x"00001021", -- addu $v0, $zero, $zero
        10 => x"00001821", -- addu $v1, $zero, $zero
        11 => x"00002021", -- addu $a0, $zero, $zero
        12 => x"00002821", -- addu $a1, $zero, $zero
        13 => x"00003021", -- addu $a2, $zero, $zero
        14 => x"00003821", -- addu $a3, $zero, $zero
        15 => x"00004021", -- addu $t0, $zero, $zero
        16 => x"00004821", -- addu $t1, $zero, $zero
        17 => x"00005021", -- addu $t2, $zero, $zero
        18 => x"00005821", -- addu $t3, $zero, $zero
        19 => x"00006021", -- addu $t4, $zero, $zero
        20 => x"00006821", -- addu $t5, $zero, $zero
        21 => x"00007021", -- addu $t6, $zero, $zero
        22 => x"00007821", -- addu $t7, $zero, $zero
        23 => x"00008021", -- addu $s0, $zero, $zero
        24 => x"00008821", -- addu $s1, $zero, $zero
        25 => x"00009021", -- addu $s2, $zero, $zero
        26 => x"00009821", -- addu $s3, $zero, $zero
        27 => x"0000A021", -- addu $s4, $zero, $zero
        28 => x"0000A821", -- addu $s5, $zero, $zero
        29 => x"0000B021", -- addu $s6, $zero, $zero
        30 => x"0000B821", -- addu $s7, $zero, $zero
        31 => x"0000C021", -- addu $t8, $zero, $zero
        32 => x"0000C821", -- addu $t9, $zero, $zero
        33 => x"0000D021", -- addu $k0, $zero, $zero
        34 => x"0000D821", -- addu $k1, $zero, $zero
        35 => x"0000E021", -- addu $gp, $zero, $zero
        36 => x"0000F821", -- addu $ra, $zero, $zero
        37 => x"3C1D0000", -- lui $sp, 0000
        38 => x"27BD0FF8", -- addiu $sp, $sp, 4088
        39 => x"0C0000F7", -- jal 247
        40 => x"03A0F021", -- addu $fp, $sp, $zero
        41 => x"08000029", -- j 41
        42 => x"00000000", -- nop
        43 => x"10C00006", -- beq $a2, $zero, 6
        44 => x"30A500FF", -- andi $a1, $a1, 00ff
        45 => x"00001021", -- addu $v0, $zero, $zero
        46 => x"24420001", -- addiu $v0, $v0, 1
        47 => x"A0850000", -- sb $a1, 0(a0)
        48 => x"1446FFFD", -- bne $v0, $a2, -3
        49 => x"24840001", -- addiu $a0, $a0, 1
        50 => x"03E00008", -- jr $ra
        51 => x"00000000", -- nop
        52 => x"04800003", -- bltz $a0, 3
        53 => x"00801021", -- addu $v0, $a0, $zero
        54 => x"03E00008", -- jr $ra
        55 => x"00000000", -- nop
        56 => x"03E00008", -- jr $ra
        57 => x"00041023", -- subu $v0, $zero, $a0
        58 => x"8F820850", -- lw $v0, 2128(gp)
        59 => x"27BDFFC8", -- addiu $sp, $sp, -56
        60 => x"00A2102A", -- slt $v0, $a1, $v0
        61 => x"AFBF0034", -- sw $ra, 52(sp)
        62 => x"AFBE0030", -- sw $fp, 48(sp)
        63 => x"AFB7002C", -- sw $s7, 44(sp)
        64 => x"AFB60028", -- sw $s6, 40(sp)
        65 => x"AFB50024", -- sw $s5, 36(sp)
        66 => x"AFB40020", -- sw $s4, 32(sp)
        67 => x"AFB3001C", -- sw $s3, 28(sp)
        68 => x"AFB20018", -- sw $s2, 24(sp)
        69 => x"AFB10014", -- sw $s1, 20(sp)
        70 => x"AFB00010", -- sw $s0, 16(sp)
        71 => x"AFA5003C", -- sw $a1, 60(sp)
        72 => x"10400039", -- beq $v0, $zero, 57
        73 => x"AFA40038", -- sw $a0, 56(sp)
        74 => x"8F85084C", -- lw $a1, 2124(gp)
        75 => x"00000000", -- nop
        76 => x"1085006D", -- beq $a0, $a1, 109
        77 => x"0000B021", -- addu $s6, $zero, $zero
        78 => x"241E0001", -- addiu $fp, $zero, 1
        79 => x"24970001", -- addiu $s7, $a0, 1
        80 => x"00161940", -- sll $v1, $s6, 10
        81 => x"001610C0", -- sll $v0, $s6, 6
        82 => x"00431021", -- addu $v0, $v0, $v1
        83 => x"3C030000", -- lui $v1, 0000
        84 => x"246308B0", -- addiu $v1, $v1, 2224
        85 => x"0062A021", -- addu $s4, $v1, $v0
        86 => x"0000A821", -- addu $s5, $zero, $zero
        87 => x"8FA30038", -- lw $v1, 56(sp)
        88 => x"00000000", -- nop
        89 => x"10600034", -- beq $v1, $zero, 52
        90 => x"00000000", -- nop
        91 => x"8E820000", -- lw $v0, 0(s4)
        92 => x"00000000", -- nop
        93 => x"1440001D", -- bne $v0, $zero, 29
        94 => x"00000000", -- nop
        95 => x"12C00005", -- beq $s6, $zero, 5
        96 => x"00001821", -- addu $v1, $zero, $zero
        97 => x"8E82FFD8", -- lw $v0, -40(s4)
        98 => x"00000000", -- nop
        99 => x"38420001", -- xori $v0, $v0, 0001
       100 => x"2C430001", -- sltiu $v1, $v0, 1
       101 => x"12A00006", -- beq $s5, $zero, 6
       102 => x"24020004", -- addiu $v0, $zero, 4
       103 => x"8E82FFFC", -- lw $v0, -4(s4)
       104 => x"00000000", -- nop
       105 => x"105E004C", -- beq $v0, $fp, 76
       106 => x"00000000", -- nop
       107 => x"24020004", -- addiu $v0, $zero, 4
       108 => x"12C20006", -- beq $s6, $v0, 6
       109 => x"24020004", -- addiu $v0, $zero, 4
       110 => x"8E820028", -- lw $v0, 40(s4)
       111 => x"00000000", -- nop
       112 => x"105E0047", -- beq $v0, $fp, 71
       113 => x"00000000", -- nop
       114 => x"24020004", -- addiu $v0, $zero, 4
       115 => x"12A20005", -- beq $s5, $v0, 5
       116 => x"00000000", -- nop
       117 => x"8E820004", -- lw $v0, 4(s4)
       118 => x"00000000", -- nop
       119 => x"105E0016", -- beq $v0, $fp, 22
       120 => x"00000000", -- nop
       121 => x"14600014", -- bne $v1, $zero, 20
       122 => x"00000000", -- nop
       123 => x"26B50001", -- addiu $s5, $s5, 1
       124 => x"24020005", -- addiu $v0, $zero, 5
       125 => x"16A2FFD9", -- bne $s5, $v0, -39
       126 => x"26940004", -- addiu $s4, $s4, 4
       127 => x"26D60001", -- addiu $s6, $s6, 1
       128 => x"16C2FFD0", -- bne $s6, $v0, -48
       129 => x"00161940", -- sll $v1, $s6, 10
       130 => x"8FBF0034", -- lw $ra, 52(sp)
       131 => x"8FBE0030", -- lw $fp, 48(sp)
       132 => x"8FB7002C", -- lw $s7, 44(sp)
       133 => x"8FB60028", -- lw $s6, 40(sp)
       134 => x"8FB50024", -- lw $s5, 36(sp)
       135 => x"8FB40020", -- lw $s4, 32(sp)
       136 => x"8FB3001C", -- lw $s3, 28(sp)
       137 => x"8FB20018", -- lw $s2, 24(sp)
       138 => x"8FB10014", -- lw $s1, 20(sp)
       139 => x"8FB00010", -- lw $s0, 16(sp)
       140 => x"03E00008", -- jr $ra
       141 => x"27BD0038", -- addiu $sp, $sp, 56
       142 => x"18A00025", -- blez $a1, 37
       143 => x"AE9E0000", -- sw $fp, 0(s4)
       144 => x"3C100000", -- lui $s0, 0000
       145 => x"3C130000", -- lui $s3, 0000
       146 => x"3C120000", -- lui $s2, 0000
       147 => x"26100A40", -- addiu $s0, $s0, 2624
       148 => x"26730854", -- addiu $s3, $s3, 2132
       149 => x"26520888", -- addiu $s2, $s2, 2184
       150 => x"080000A4", -- j 164
       151 => x"00008821", -- addu $s1, $zero, $zero
       152 => x"8FA5003C", -- lw $a1, 60(sp)
       153 => x"04400018", -- bltz $v0, 24
       154 => x"00651821", -- addu $v1, $v1, $a1
       155 => x"0C00003A", -- jal 58
       156 => x"00622821", -- addu $a1, $v1, $v0
       157 => x"8F85084C", -- lw $a1, 2124(gp)
       158 => x"AE000000", -- sw $zero, 0(s0)
       159 => x"0225102A", -- slt $v0, $s1, $a1
       160 => x"26100004", -- addiu $s0, $s0, 4
       161 => x"26730004", -- addiu $s3, $s3, 4
       162 => x"10400011", -- beq $v0, $zero, 17
       163 => x"26520004", -- addiu $s2, $s2, 4
       164 => x"8E020000", -- lw $v0, 0(s0)
       165 => x"26310001", -- addiu $s1, $s1, 1
       166 => x"1440FFF8", -- bne $v0, $zero, -8
       167 => x"02E02021", -- addu $a0, $s7, $zero
       168 => x"8E630000", -- lw $v1, 0(s3)
       169 => x"8E420000", -- lw $v0, 0(s2)
       170 => x"00761823", -- subu $v1, $v1, $s6
       171 => x"AE1E0000", -- sw $fp, 0(s0)
       172 => x"0461FFEB", -- bgez $v1, -21
       173 => x"00551023", -- subu $v0, $v0, $s5
       174 => x"8FA5003C", -- lw $a1, 60(sp)
       175 => x"00031823", -- subu $v1, $zero, $v1
       176 => x"0441FFEA", -- bgez $v0, -22
       177 => x"00651821", -- addu $v1, $v1, $a1
       178 => x"0800009B", -- j 155
       179 => x"00021023", -- subu $v0, $zero, $v0
       180 => x"0800007B", -- j 123
       181 => x"AE800000", -- sw $zero, 0(s4)
       182 => x"0800006B", -- j 107
       183 => x"24030001", -- addiu $v1, $zero, 1
       184 => x"08000072", -- j 114
       185 => x"24030001", -- addiu $v1, $zero, 1
       186 => x"8FA2003C", -- lw $v0, 60(sp)
       187 => x"08000082", -- j 130
       188 => x"AF820850", -- sw $v0, 2128(gp)
       189 => x"27BDFFE8", -- addiu $sp, $sp, -24
       190 => x"3C020000", -- lui $v0, 0000
       191 => x"3C030000", -- lui $v1, 0000
       192 => x"AFBF0014", -- sw $ra, 20(sp)
       193 => x"AF80084C", -- sw $zero, 2124(gp)
       194 => x"00803021", -- addu $a2, $a0, $zero
       195 => x"244A0854", -- addiu $t2, $v0, 2132
       196 => x"246B0888", -- addiu $t3, $v1, 2184
       197 => x"00003821", -- addu $a3, $zero, $zero
       198 => x"2409002A", -- addiu $t1, $zero, 42
       199 => x"24080005", -- addiu $t0, $zero, 5
       200 => x"00002821", -- addu $a1, $zero, $zero
       201 => x"00C51021", -- addu $v0, $a2, $a1
       202 => x"80430000", -- lb $v1, 0(v0)
       203 => x"00000000", -- nop
       204 => x"10690020", -- beq $v1, $t1, 32
       205 => x"00000000", -- nop
       206 => x"24A50001", -- addiu $a1, $a1, 1
       207 => x"14A8FFFA", -- bne $a1, $t0, -6
       208 => x"00C51021", -- addu $v0, $a2, $a1
       209 => x"24E70001", -- addiu $a3, $a3, 1
       210 => x"14E5FFF5", -- bne $a3, $a1, -11
       211 => x"24C60005", -- addiu $a2, $a2, 5
       212 => x"3C020000", -- lui $v0, 0000
       213 => x"3C030000", -- lui $v1, 0000
       214 => x"244208B0", -- addiu $v0, $v0, 2224
       215 => x"24630A40", -- addiu $v1, $v1, 2624
       216 => x"A0400000", -- sb $zero, 0(v0)
       217 => x"24420001", -- addiu $v0, $v0, 1
       218 => x"1443FFFD", -- bne $v0, $v1, -3
       219 => x"00000000", -- nop
       220 => x"3C020000", -- lui $v0, 0000
       221 => x"3C030000", -- lui $v1, 0000
       222 => x"24420A40", -- addiu $v0, $v0, 2624
       223 => x"24630A68", -- addiu $v1, $v1, 2664
       224 => x"A0400000", -- sb $zero, 0(v0)
       225 => x"24420001", -- addiu $v0, $v0, 1
       226 => x"1443FFFD", -- bne $v0, $v1, -3
       227 => x"00002021", -- addu $a0, $zero, $zero
       228 => x"3C02000F", -- lui $v0, 000f
       229 => x"34424240", -- ori $v0, $v0, 4240
       230 => x"00002821", -- addu $a1, $zero, $zero
       231 => x"0C00003A", -- jal 58
       232 => x"AF820850", -- sw $v0, 2128(gp)
       233 => x"8FBF0014", -- lw $ra, 20(sp)
       234 => x"8F820850", -- lw $v0, 2128(gp)
       235 => x"03E00008", -- jr $ra
       236 => x"27BD0018", -- addiu $sp, $sp, 24
       237 => x"8F82084C", -- lw $v0, 2124(gp)
       238 => x"00000000", -- nop
       239 => x"00021880", -- sll $v1, $v0, 4
       240 => x"006B2021", -- addu $a0, $v1, $t3
       241 => x"24420001", -- addiu $v0, $v0, 1
       242 => x"006A1821", -- addu $v1, $v1, $t2
       243 => x"AC850000", -- sw $a1, 0(a0)
       244 => x"AC670000", -- sw $a3, 0(v1)
       245 => x"080000CE", -- j 206
       246 => x"AF82084C", -- sw $v0, 2124(gp)
       247 => x"27BDFFE0", -- addiu $sp, $sp, -32
       248 => x"3C020000", -- lui $v0, 0000
       249 => x"AFB00010", -- sw $s0, 16(sp)
       250 => x"3C030000", -- lui $v1, 0000
       251 => x"24500800", -- addiu $s0, $v0, 2048
       252 => x"3C020000", -- lui $v0, 0000
       253 => x"AFB20018", -- sw $s2, 24(sp)
       254 => x"AFB10014", -- sw $s1, 20(sp)
       255 => x"AFBF001C", -- sw $ra, 28(sp)
       256 => x"2471087C", -- addiu $s1, $v1, 2172
       257 => x"2452084B", -- addiu $s2, $v0, 2123
       258 => x"0C0000BD", -- jal 189
       259 => x"02002021", -- addu $a0, $s0, $zero
       260 => x"26100019", -- addiu $s0, $s0, 25
       261 => x"AE220000", -- sw $v0, 0(s1)
       262 => x"1650FFFB", -- bne $s2, $s0, -5
       263 => x"26310004", -- addiu $s1, $s1, 4
       264 => x"8FBF001C", -- lw $ra, 28(sp)
       265 => x"00001021", -- addu $v0, $zero, $zero
       266 => x"8FB20018", -- lw $s2, 24(sp)
       267 => x"8FB10014", -- lw $s1, 20(sp)
       268 => x"8FB00010", -- lw $s0, 16(sp)
       269 => x"03E00008", -- jr $ra
       270 => x"27BD0020", -- addiu $sp, $sp, 32
       271 => x"00000000", -- nop
       272 => x"00000000", -- nop
       273 => x"00000000", -- nop
       274 => x"00000000", -- nop
       275 => x"00000000", -- nop
       276 => x"00000000", -- nop
       277 => x"00000000", -- nop
       278 => x"00000000", -- nop
       279 => x"00000000", -- nop
       280 => x"00000000", -- nop
       281 => x"00000000", -- nop
       282 => x"00000000", -- nop
       283 => x"00000000", -- nop
       284 => x"00000000", -- nop
       285 => x"00000000", -- nop
       286 => x"00000000", -- nop
       287 => x"00000000", -- nop
       288 => x"00000000", -- nop
       289 => x"00000000", -- nop
       290 => x"00000000", -- nop
       291 => x"00000000", -- nop
       292 => x"00000000", -- nop
       293 => x"00000000", -- nop
       294 => x"00000000", -- nop
       295 => x"00000000", -- nop
       296 => x"00000000", -- nop
       297 => x"00000000", -- nop
       298 => x"00000000", -- nop
       299 => x"00000000", -- nop
       300 => x"00000000", -- nop
       301 => x"00000000", -- nop
       302 => x"00000000", -- nop
       303 => x"00000000", -- nop
       304 => x"00000000", -- nop
       305 => x"00000000", -- nop
       306 => x"00000000", -- nop
       307 => x"00000000", -- nop
       308 => x"00000000", -- nop
       309 => x"00000000", -- nop
       310 => x"00000000", -- nop
       311 => x"00000000", -- nop
       312 => x"00000000", -- nop
       313 => x"00000000", -- nop
       314 => x"00000000", -- nop
       315 => x"00000000", -- nop
       316 => x"00000000", -- nop
       317 => x"00000000", -- nop
       318 => x"00000000", -- nop
       319 => x"00000000", -- nop
       320 => x"00000000", -- nop
       321 => x"00000000", -- nop
       322 => x"00000000", -- nop
       323 => x"00000000", -- nop
       324 => x"00000000", -- nop
       325 => x"00000000", -- nop
       326 => x"00000000", -- nop
       327 => x"00000000", -- nop
       328 => x"00000000", -- nop
       329 => x"00000000", -- nop
       330 => x"00000000", -- nop
       331 => x"00000000", -- nop
       332 => x"00000000", -- nop
       333 => x"00000000", -- nop
       334 => x"00000000", -- nop
       335 => x"00000000", -- nop
       336 => x"00000000", -- nop
       337 => x"00000000", -- nop
       338 => x"00000000", -- nop
       339 => x"00000000", -- nop
       340 => x"00000000", -- nop
       341 => x"00000000", -- nop
       342 => x"00000000", -- nop
       343 => x"00000000", -- nop
       344 => x"00000000", -- nop
       345 => x"00000000", -- nop
       346 => x"00000000", -- nop
       347 => x"00000000", -- nop
       348 => x"00000000", -- nop
       349 => x"00000000", -- nop
       350 => x"00000000", -- nop
       351 => x"00000000", -- nop
       352 => x"00000000", -- nop
       353 => x"00000000", -- nop
       354 => x"00000000", -- nop
       355 => x"00000000", -- nop
       356 => x"00000000", -- nop
       357 => x"00000000", -- nop
       358 => x"00000000", -- nop
       359 => x"00000000", -- nop
       360 => x"00000000", -- nop
       361 => x"00000000", -- nop
       362 => x"00000000", -- nop
       363 => x"00000000", -- nop
       364 => x"00000000", -- nop
       365 => x"00000000", -- nop
       366 => x"00000000", -- nop
       367 => x"00000000", -- nop
       368 => x"00000000", -- nop
       369 => x"00000000", -- nop
       370 => x"00000000", -- nop
       371 => x"00000000", -- nop
       372 => x"00000000", -- nop
       373 => x"00000000", -- nop
       374 => x"00000000", -- nop
       375 => x"00000000", -- nop
       376 => x"00000000", -- nop
       377 => x"00000000", -- nop
       378 => x"00000000", -- nop
       379 => x"00000000", -- nop
       380 => x"00000000", -- nop
       381 => x"00000000", -- nop
       382 => x"00000000", -- nop
       383 => x"00000000", -- nop
       384 => x"00000000", -- nop
       385 => x"00000000", -- nop
       386 => x"00000000", -- nop
       387 => x"00000000", -- nop
       388 => x"00000000", -- nop
       389 => x"00000000", -- nop
       390 => x"00000000", -- nop
       391 => x"00000000", -- nop
       392 => x"00000000", -- nop
       393 => x"00000000", -- nop
       394 => x"00000000", -- nop
       395 => x"00000000", -- nop
       396 => x"00000000", -- nop
       397 => x"00000000", -- nop
       398 => x"00000000", -- nop
       399 => x"00000000", -- nop
       400 => x"00000000", -- nop
       401 => x"00000000", -- nop
       402 => x"00000000", -- nop
       403 => x"00000000", -- nop
       404 => x"00000000", -- nop
       405 => x"00000000", -- nop
       406 => x"00000000", -- nop
       407 => x"00000000", -- nop
       408 => x"00000000", -- nop
       409 => x"00000000", -- nop
       410 => x"00000000", -- nop
       411 => x"00000000", -- nop
       412 => x"00000000", -- nop
       413 => x"00000000", -- nop
       414 => x"00000000", -- nop
       415 => x"00000000", -- nop
       416 => x"00000000", -- nop
       417 => x"00000000", -- nop
       418 => x"00000000", -- nop
       419 => x"00000000", -- nop
       420 => x"00000000", -- nop
       421 => x"00000000", -- nop
       422 => x"00000000", -- nop
       423 => x"00000000", -- nop
       424 => x"00000000", -- nop
       425 => x"00000000", -- nop
       426 => x"00000000", -- nop
       427 => x"00000000", -- nop
       428 => x"00000000", -- nop
       429 => x"00000000", -- nop
       430 => x"00000000", -- nop
       431 => x"00000000", -- nop
       432 => x"00000000", -- nop
       433 => x"00000000", -- nop
       434 => x"00000000", -- nop
       435 => x"00000000", -- nop
       436 => x"00000000", -- nop
       437 => x"00000000", -- nop
       438 => x"00000000", -- nop
       439 => x"00000000", -- nop
       440 => x"00000000", -- nop
       441 => x"00000000", -- nop
       442 => x"00000000", -- nop
       443 => x"00000000", -- nop
       444 => x"00000000", -- nop
       445 => x"00000000", -- nop
       446 => x"00000000", -- nop
       447 => x"00000000", -- nop
       448 => x"00000000", -- nop
       449 => x"00000000", -- nop
       450 => x"00000000", -- nop
       451 => x"00000000", -- nop
       452 => x"00000000", -- nop
       453 => x"00000000", -- nop
       454 => x"00000000", -- nop
       455 => x"00000000", -- nop
       456 => x"00000000", -- nop
       457 => x"00000000", -- nop
       458 => x"00000000", -- nop
       459 => x"00000000", -- nop
       460 => x"00000000", -- nop
       461 => x"00000000", -- nop
       462 => x"00000000", -- nop
       463 => x"00000000", -- nop
       464 => x"00000000", -- nop
       465 => x"00000000", -- nop
       466 => x"00000000", -- nop
       467 => x"00000000", -- nop
       468 => x"00000000", -- nop
       469 => x"00000000", -- nop
       470 => x"00000000", -- nop
       471 => x"00000000", -- nop
       472 => x"00000000", -- nop
       473 => x"00000000", -- nop
       474 => x"00000000", -- nop
       475 => x"00000000", -- nop
       476 => x"00000000", -- nop
       477 => x"00000000", -- nop
       478 => x"00000000", -- nop
       479 => x"00000000", -- nop
       480 => x"00000000", -- nop
       481 => x"00000000", -- nop
       482 => x"00000000", -- nop
       483 => x"00000000", -- nop
       484 => x"00000000", -- nop
       485 => x"00000000", -- nop
       486 => x"00000000", -- nop
       487 => x"00000000", -- nop
       488 => x"00000000", -- nop
       489 => x"00000000", -- nop
       490 => x"00000000", -- nop
       491 => x"00000000", -- nop
       492 => x"00000000", -- nop
       493 => x"00000000", -- nop
       494 => x"00000000", -- nop
       495 => x"00000000", -- nop
       496 => x"00000000", -- nop
       497 => x"00000000", -- nop
       498 => x"00000000", -- nop
       499 => x"00000000", -- nop
       500 => x"00000000", -- nop
       501 => x"00000000", -- nop
       502 => x"00000000", -- nop
       503 => x"00000000", -- nop
       504 => x"00000000", -- nop
       505 => x"00000000", -- nop
       506 => x"00000000", -- nop
       507 => x"00000000", -- nop
       508 => x"00000000", -- nop
       509 => x"00000000", -- nop
       510 => x"00000000", -- nop
       511 => x"00000000"  -- nop
    );

BEGIN

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF R='1' THEN
                DATA_OUT <= TMP_RAM(CONV_INTEGER(UNSIGNED(RADDR(ADDR-1 DOWNTO 2))));
            ELSE
                DATA_OUT <= (DATA_OUT'RANGE => 'Z');
            END IF;
        END IF;
    END IF;
    END PROCESS;

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF W='1' THEN
                TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2)))) <= DATA_IN;
            END IF;
        END IF;
    END IF;
    END PROCESS;

END BEHAV_CODE;

ARCHITECTURE BEHAV_DATA OF SRAM IS

    TYPE RAM_TYPE IS ARRAY (0 TO DEPTH-1) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL IBYTE0:     STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL IBYTE1:     STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL IBYTE2:     STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL IBYTE3:     STD_LOGIC_VECTOR(7 DOWNTO 0);

    SIGNAL OBYTE:      STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL OHALF:      STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SBYTE:      STD_LOGIC_VECTOR(23 DOWNTO 0);
    SIGNAL SHALF:      STD_LOGIC_VECTOR(15 DOWNTO 0);

    SIGNAL RWORD:      STD_LOGIC_VECTOR(31 DOWNTO 0):= x"00000000";

    SIGNAL RADDR2:     STD_LOGIC_VECTOR(1 DOWNTO 0):= "00";
    SIGNAL MODE2:      STD_LOGIC_VECTOR(2 DOWNTO 0):= "000";
    SIGNAL ISSIGNED2:  STD_LOGIC:= '0';

    SIGNAL W0:         STD_LOGIC;
    SIGNAL W1:         STD_LOGIC;
    SIGNAL W2:         STD_LOGIC;
    SIGNAL W3:         STD_LOGIC;

    SIGNAL TMP_RAM: RAM_TYPE := (

         0 => x"2E2E2E2E",
         1 => x"2E2E2E2A",
         2 => x"2A2E2E2E",
         3 => x"2E2E2E2E",
         4 => x"2E2E2A2E",
         5 => x"2E2E2E2E",
         6 => x"2E2E2E2E",
         7 => x"2E2E2E2E",
         8 => x"2E2E2E2E",
         9 => x"2A2A2E2E",
        10 => x"2E2A2E2E",
        11 => x"2E2A2A2E",
        12 => x"2E2E2A2E",
        13 => x"2E2E2A2E",
        14 => x"2E2E2E2E",
        15 => x"2E2E2E2E",
        16 => x"2E2E2E2E",
        17 => x"2E2E2A2E",
        18 => x"2E2E2A00",
        19 => x"55555555",
        20 => x"55555555",
        21 => x"55555555",
        22 => x"55555555",
        23 => x"55555555",
        24 => x"55555555",
        25 => x"55555555",
        26 => x"55555555",
        27 => x"55555555",
        28 => x"55555555",
        29 => x"55555555",
        30 => x"55555555",
        31 => x"55555555",
        32 => x"55555555",
        33 => x"55555555",
        34 => x"55555555",
        35 => x"55555555",
        36 => x"55555555",
        37 => x"55555555",
        38 => x"55555555",
        39 => x"55555555",
        40 => x"55555555",
        41 => x"55555555",
        42 => x"55555555",
        43 => x"55555555",
        44 => x"55555555",
        45 => x"55555555",
        46 => x"55555555",
        47 => x"55555555",
        48 => x"55555555",
        49 => x"55555555",
        50 => x"55555555",
        51 => x"55555555",
        52 => x"55555555",
        53 => x"55555555",
        54 => x"55555555",
        55 => x"55555555",
        56 => x"55555555",
        57 => x"55555555",
        58 => x"55555555",
        59 => x"55555555",
        60 => x"55555555",
        61 => x"55555555",
        62 => x"55555555",
        63 => x"55555555",
        64 => x"55555555",
        65 => x"55555555",
        66 => x"55555555",
        67 => x"55555555",
        68 => x"55555555",
        69 => x"55555555",
        70 => x"55555555",
        71 => x"55555555",
        72 => x"55555555",
        73 => x"55555555",
        74 => x"55555555",
        75 => x"55555555",
        76 => x"55555555",
        77 => x"55555555",
        78 => x"55555555",
        79 => x"55555555",
        80 => x"55555555",
        81 => x"55555555",
        82 => x"55555555",
        83 => x"55555555",
        84 => x"55555555",
        85 => x"55555555",
        86 => x"55555555",
        87 => x"55555555",
        88 => x"55555555",
        89 => x"55555555",
        90 => x"55555555",
        91 => x"55555555",
        92 => x"55555555",
        93 => x"55555555",
        94 => x"55555555",
        95 => x"55555555",
        96 => x"55555555",
        97 => x"55555555",
        98 => x"55555555",
        99 => x"55555555",
       100 => x"55555555",
       101 => x"55555555",
       102 => x"55555555",
       103 => x"55555555",
       104 => x"55555555",
       105 => x"55555555",
       106 => x"55555555",
       107 => x"55555555",
       108 => x"55555555",
       109 => x"55555555",
       110 => x"55555555",
       111 => x"55555555",
       112 => x"55555555",
       113 => x"55555555",
       114 => x"55555555",
       115 => x"55555555",
       116 => x"55555555",
       117 => x"55555555",
       118 => x"55555555",
       119 => x"55555555",
       120 => x"55555555",
       121 => x"55555555",
       122 => x"55555555",
       123 => x"55555555",
       124 => x"55555555",
       125 => x"55555555",
       126 => x"55555555",
       127 => x"55555555",
       128 => x"55555555",
       129 => x"55555555",
       130 => x"55555555",
       131 => x"55555555",
       132 => x"55555555",
       133 => x"55555555",
       134 => x"55555555",
       135 => x"55555555",
       136 => x"55555555",
       137 => x"55555555",
       138 => x"55555555",
       139 => x"55555555",
       140 => x"55555555",
       141 => x"55555555",
       142 => x"55555555",
       143 => x"55555555",
       144 => x"55555555",
       145 => x"55555555",
       146 => x"55555555",
       147 => x"55555555",
       148 => x"55555555",
       149 => x"55555555",
       150 => x"55555555",
       151 => x"55555555",
       152 => x"55555555",
       153 => x"55555555",
       154 => x"55555555",
       155 => x"55555555",
       156 => x"55555555",
       157 => x"55555555",
       158 => x"55555555",
       159 => x"55555555",
       160 => x"55555555",
       161 => x"55555555",
       162 => x"55555555",
       163 => x"55555555",
       164 => x"55555555",
       165 => x"55555555",
       166 => x"55555555",
       167 => x"55555555",
       168 => x"55555555",
       169 => x"55555555",
       170 => x"55555555",
       171 => x"55555555",
       172 => x"55555555",
       173 => x"55555555",
       174 => x"55555555",
       175 => x"55555555",
       176 => x"55555555",
       177 => x"55555555",
       178 => x"55555555",
       179 => x"55555555",
       180 => x"55555555",
       181 => x"55555555",
       182 => x"55555555",
       183 => x"55555555",
       184 => x"55555555",
       185 => x"55555555",
       186 => x"55555555",
       187 => x"55555555",
       188 => x"55555555",
       189 => x"55555555",
       190 => x"55555555",
       191 => x"55555555",
       192 => x"55555555",
       193 => x"55555555",
       194 => x"55555555",
       195 => x"55555555",
       196 => x"55555555",
       197 => x"55555555",
       198 => x"55555555",
       199 => x"55555555",
       200 => x"55555555",
       201 => x"55555555",
       202 => x"55555555",
       203 => x"55555555",
       204 => x"55555555",
       205 => x"55555555",
       206 => x"55555555",
       207 => x"55555555",
       208 => x"55555555",
       209 => x"55555555",
       210 => x"55555555",
       211 => x"55555555",
       212 => x"55555555",
       213 => x"55555555",
       214 => x"55555555",
       215 => x"55555555",
       216 => x"55555555",
       217 => x"55555555",
       218 => x"55555555",
       219 => x"55555555",
       220 => x"55555555",
       221 => x"55555555",
       222 => x"55555555",
       223 => x"55555555",
       224 => x"55555555",
       225 => x"55555555",
       226 => x"55555555",
       227 => x"55555555",
       228 => x"55555555",
       229 => x"55555555",
       230 => x"55555555",
       231 => x"55555555",
       232 => x"55555555",
       233 => x"55555555",
       234 => x"55555555",
       235 => x"55555555",
       236 => x"55555555",
       237 => x"55555555",
       238 => x"55555555",
       239 => x"55555555",
       240 => x"55555555",
       241 => x"55555555",
       242 => x"55555555",
       243 => x"55555555",
       244 => x"55555555",
       245 => x"55555555",
       246 => x"55555555",
       247 => x"55555555",
       248 => x"55555555",
       249 => x"55555555",
       250 => x"55555555",
       251 => x"55555555",
       252 => x"55555555",
       253 => x"55555555",
       254 => x"55555555",
       255 => x"55555555",
       256 => x"55555555",
       257 => x"55555555",
       258 => x"55555555",
       259 => x"55555555",
       260 => x"55555555",
       261 => x"55555555",
       262 => x"55555555",
       263 => x"55555555",
       264 => x"55555555",
       265 => x"55555555",
       266 => x"55555555",
       267 => x"55555555",
       268 => x"55555555",
       269 => x"55555555",
       270 => x"55555555",
       271 => x"55555555",
       272 => x"55555555",
       273 => x"55555555",
       274 => x"55555555",
       275 => x"55555555",
       276 => x"55555555",
       277 => x"55555555",
       278 => x"55555555",
       279 => x"55555555",
       280 => x"55555555",
       281 => x"55555555",
       282 => x"55555555",
       283 => x"55555555",
       284 => x"55555555",
       285 => x"55555555",
       286 => x"55555555",
       287 => x"55555555",
       288 => x"55555555",
       289 => x"55555555",
       290 => x"55555555",
       291 => x"55555555",
       292 => x"55555555",
       293 => x"55555555",
       294 => x"55555555",
       295 => x"55555555",
       296 => x"55555555",
       297 => x"55555555",
       298 => x"55555555",
       299 => x"55555555",
       300 => x"55555555",
       301 => x"55555555",
       302 => x"55555555",
       303 => x"55555555",
       304 => x"55555555",
       305 => x"55555555",
       306 => x"55555555",
       307 => x"55555555",
       308 => x"55555555",
       309 => x"55555555",
       310 => x"55555555",
       311 => x"55555555",
       312 => x"55555555",
       313 => x"55555555",
       314 => x"55555555",
       315 => x"55555555",
       316 => x"55555555",
       317 => x"55555555",
       318 => x"55555555",
       319 => x"55555555",
       320 => x"55555555",
       321 => x"55555555",
       322 => x"55555555",
       323 => x"55555555",
       324 => x"55555555",
       325 => x"55555555",
       326 => x"55555555",
       327 => x"55555555",
       328 => x"55555555",
       329 => x"55555555",
       330 => x"55555555",
       331 => x"55555555",
       332 => x"55555555",
       333 => x"55555555",
       334 => x"55555555",
       335 => x"55555555",
       336 => x"55555555",
       337 => x"55555555",
       338 => x"55555555",
       339 => x"55555555",
       340 => x"55555555",
       341 => x"55555555",
       342 => x"55555555",
       343 => x"55555555",
       344 => x"55555555",
       345 => x"55555555",
       346 => x"55555555",
       347 => x"55555555",
       348 => x"55555555",
       349 => x"55555555",
       350 => x"55555555",
       351 => x"55555555",
       352 => x"55555555",
       353 => x"55555555",
       354 => x"55555555",
       355 => x"55555555",
       356 => x"55555555",
       357 => x"55555555",
       358 => x"55555555",
       359 => x"55555555",
       360 => x"55555555",
       361 => x"55555555",
       362 => x"55555555",
       363 => x"55555555",
       364 => x"55555555",
       365 => x"55555555",
       366 => x"55555555",
       367 => x"55555555",
       368 => x"55555555",
       369 => x"55555555",
       370 => x"55555555",
       371 => x"55555555",
       372 => x"55555555",
       373 => x"55555555",
       374 => x"55555555",
       375 => x"55555555",
       376 => x"55555555",
       377 => x"55555555",
       378 => x"55555555",
       379 => x"55555555",
       380 => x"55555555",
       381 => x"55555555",
       382 => x"55555555",
       383 => x"55555555",
       384 => x"55555555",
       385 => x"55555555",
       386 => x"55555555",
       387 => x"55555555",
       388 => x"55555555",
       389 => x"55555555",
       390 => x"55555555",
       391 => x"55555555",
       392 => x"55555555",
       393 => x"55555555",
       394 => x"55555555",
       395 => x"55555555",
       396 => x"55555555",
       397 => x"55555555",
       398 => x"55555555",
       399 => x"55555555",
       400 => x"55555555",
       401 => x"55555555",
       402 => x"55555555",
       403 => x"55555555",
       404 => x"55555555",
       405 => x"55555555",
       406 => x"55555555",
       407 => x"55555555",
       408 => x"55555555",
       409 => x"55555555",
       410 => x"55555555",
       411 => x"55555555",
       412 => x"55555555",
       413 => x"55555555",
       414 => x"55555555",
       415 => x"55555555",
       416 => x"55555555",
       417 => x"55555555",
       418 => x"55555555",
       419 => x"55555555",
       420 => x"55555555",
       421 => x"55555555",
       422 => x"55555555",
       423 => x"55555555",
       424 => x"55555555",
       425 => x"55555555",
       426 => x"55555555",
       427 => x"55555555",
       428 => x"55555555",
       429 => x"55555555",
       430 => x"55555555",
       431 => x"55555555",
       432 => x"55555555",
       433 => x"55555555",
       434 => x"55555555",
       435 => x"55555555",
       436 => x"55555555",
       437 => x"55555555",
       438 => x"55555555",
       439 => x"55555555",
       440 => x"55555555",
       441 => x"55555555",
       442 => x"55555555",
       443 => x"55555555",
       444 => x"55555555",
       445 => x"55555555",
       446 => x"55555555",
       447 => x"55555555",
       448 => x"55555555",
       449 => x"55555555",
       450 => x"55555555",
       451 => x"55555555",
       452 => x"55555555",
       453 => x"55555555",
       454 => x"55555555",
       455 => x"55555555",
       456 => x"55555555",
       457 => x"55555555",
       458 => x"55555555",
       459 => x"55555555",
       460 => x"55555555",
       461 => x"55555555",
       462 => x"55555555",
       463 => x"55555555",
       464 => x"55555555",
       465 => x"55555555",
       466 => x"55555555",
       467 => x"55555555",
       468 => x"55555555",
       469 => x"55555555",
       470 => x"55555555",
       471 => x"55555555",
       472 => x"55555555",
       473 => x"55555555",
       474 => x"55555555",
       475 => x"55555555",
       476 => x"55555555",
       477 => x"55555555",
       478 => x"55555555",
       479 => x"55555555",
       480 => x"55555555",
       481 => x"55555555",
       482 => x"55555555",
       483 => x"55555555",
       484 => x"55555555",
       485 => x"55555555",
       486 => x"55555555",
       487 => x"55555555",
       488 => x"55555555",
       489 => x"55555555",
       490 => x"55555555",
       491 => x"55555555",
       492 => x"55555555",
       493 => x"55555555",
       494 => x"55555555",
       495 => x"55555555",
       496 => x"55555555",
       497 => x"55555555",
       498 => x"55555555",
       499 => x"55555555",
       500 => x"55555555",
       501 => x"55555555",
       502 => x"55555555",
       503 => x"55555555",
       504 => x"55555555",
       505 => x"55555555",
       506 => x"55555555",
       507 => x"55555555",
       508 => x"55555555",
       509 => x"55555555",
       510 => x"55555555",
       511 => x"55555555"
    );

BEGIN
    -- READ LOGIC
    OBYTE    <=      RWORD(31 DOWNTO 24) WHEN RADDR2(1 DOWNTO 0) = "00"
                ELSE RWORD(23 DOWNTO 16) WHEN RADDR2(1 DOWNTO 0) = "01"
                ELSE RWORD(15 DOWNTO  8) WHEN RADDR2(1 DOWNTO 0) = "10"
                ELSE RWORD( 7 DOWNTO  0);

    OHALF    <=      RWORD(31 DOWNTO 16) WHEN RADDR2(1 DOWNTO 0) = "00"
                ELSE RWORD(15 DOWNTO  0); -- THIS IS CASE "11", WE DON'T HANDLE THE OTHER CASES


    SBYTE    <=      x"FFFFFF" WHEN (OBYTE(7)  AND ISSIGNED2) = '1' ELSE x"000000";
    SHALF    <=      x"FFFF"   WHEN (OHALF(15) AND ISSIGNED2) = '1' ELSE x"0000";


    DATA_OUT <=      SBYTE & OBYTE WHEN MODE2(2) = '1'
                ELSE SHALF & OHALF WHEN MODE2(1) = '1'
                ELSE RWORD WHEN MODE2(0) = '1';

    -- WRITE LOGIC

    IBYTE0 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN(15 DOWNTO 8) WHEN MODE(1)='1' ELSE DATA_IN(31 DOWNTO  24);
    IBYTE1 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN( 7 DOWNTO 0) WHEN MODE(1)='1' ELSE DATA_IN(23 DOWNTO  16);
    IBYTE2 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN(15 DOWNTO 8) WHEN MODE(1)='1' ELSE DATA_IN(15 DOWNTO   8);
    IBYTE3 <= DATA_IN(7 DOWNTO  0) WHEN MODE(2)='1' ELSE DATA_IN( 7 DOWNTO 0) WHEN MODE(1)='1' ELSE DATA_IN( 7 DOWNTO   0);

    W0 <= (   (MODE(2) AND NOT(WADDR(1) OR   WADDR(0)))  --B: "00"
           OR (MODE(1) AND NOT(WADDR(1)))                --H: "0x"
           OR  MODE(0)) AND W;                           --W: "Xx"
    W1 <= (   (MODE(2) AND NOT(WADDR(1)) AND WADDR(0))   --B: "01"
           OR (MODE(1) AND NOT(WADDR(1)))                --H: "0x"
           OR  MODE(0)) AND W;                           --W: "Xx"
    W2 <= (   (MODE(2) AND NOT(WADDR(0)) AND WADDR(1))   --B: "10"
           OR (MODE(1) AND     WADDR(1))                 --H: "1x"
           OR  MODE(0)) AND W;                           --W: "Xx"
    W3 <= (   (MODE(2) AND     WADDR(1) AND  WADDR(0))   --B: "11"
           OR (MODE(1) AND     WADDR(1))                 --H: "1x"
           OR  MODE(0)) AND W;                           --W: "Xx"

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        MODE2     <= MODE;
        ISSIGNED2 <= ISSIGNED;
        RADDR2 <= RADDR(1 DOWNTO 0);
    END IF;
    END PROCESS;

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF R='1' THEN
                RWORD <= TMP_RAM(CONV_INTEGER(UNSIGNED(RADDR(ADDR-1 DOWNTO 2))));
            ELSE
                RWORD <= (DATA_OUT'RANGE => 'Z');
            END IF;
        END IF;
    END IF;
    END PROCESS;

    PROCESS(CLK)
    BEGIN
    IF (CLK'EVENT AND CLK='1') THEN
        IF ENABLE='1' THEN
            IF W='1' THEN
                IF W0 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(31 DOWNTO 24) <= IBYTE0;
                END IF;
                IF W1 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(23 DOWNTO 16) <= IBYTE1;
                END IF;
                IF W2 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(15 DOWNTO  8) <= IBYTE2;
                END IF;
                IF W3 = '1' THEN
                    TMP_RAM(CONV_INTEGER(UNSIGNED(WADDR(ADDR-1 DOWNTO 2))))(7  DOWNTO  0) <= IBYTE3;
                END IF;
            END IF;
        END IF;
    END IF;
    END PROCESS;

END BEHAV_DATA;
